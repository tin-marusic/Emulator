parameter integer matrixE [0:1743] = {
/* num inputs = 138 (in0-in137) */
/* num outputs = 428(out0-out427) */
//* max inputs per outputs = 9 */
//* total number of input in adders 658 */

/* out0000_em-eta16-phi16 */     0, 
/* out0001_em-eta16-phi17 */     0, 
/* out0002_em-eta16-phi18 */     0, 
/* out0003_em-eta16-phi19 */     0, 
/* out0004_em-eta17-phi15 */     0, 
/* out0005_em-eta17-phi16 */     0, 
/* out0006_em-eta17-phi17 */     0, 
/* out0007_em-eta17-phi18 */     0, 
/* out0008_em-eta12-phi19 */     0, 
/* out0009_em-eta12-phi20 */     1, 58, 1, 
/* out0010_em-eta12-phi21 */     1, 58, 1, 
/* out0011_em-eta13-phi18 */     0, 
/* out0012_em-eta13-phi19 */     0, 
/* out0013_em-eta13-phi20 */     0, 
/* out0014_em-eta13-phi21 */     0, 
/* out0015_em-eta14-phi20 */     0, 
/* out0016_em-eta9-phi20 */     1, 93, 1, 
/* out0017_em-eta9-phi21 */     2, 59, 1, 110, 1, 
/* out0018_em-eta9-phi22 */     2, 59, 1, 110, 1, 
/* out0019_em-eta10-phi20 */     1, 58, 1, 
/* out0020_em-eta10-phi21 */     1, 58, 1, 
/* out0021_em-eta10-phi22 */     1, 58, 1, 
/* out0022_em-eta11-phi20 */     1, 58, 1, 
/* out0023_em-eta11-phi21 */     1, 58, 1, 
/* out0024_em-eta6-phi21 */     0, 
/* out0025_em-eta6-phi22 */     0, 
/* out0026_em-eta7-phi20 */     0, 
/* out0027_em-eta7-phi21 */     2, 59, 1, 110, 1, 
/* out0028_em-eta7-phi22 */     1, 59, 1, 
/* out0029_em-eta8-phi21 */     2, 59, 2, 110, 2, 
/* out0030_em-eta8-phi22 */     2, 59, 1, 110, 2, 
/* out0031_em-eta4-phi21 */     0, 
/* out0032_em-eta4-phi22 */     0, 
/* out0033_em-eta5-phi21 */     0, 
/* out0034_em-eta5-phi22 */     0, 
/* out0035_em-eta5-phi23 */     0, 
/* out0036_em-eta2-phi22 */     0, 
/* out0037_em-eta3-phi21 */     0, 
/* out0038_em-eta3-phi22 */     0, 
/* out0039_em-eta3-phi23 */     0, 
/* out0040_em-eta1-phi22 */     1, 22, 1, 
/* out0041_em-eta1-phi23 */     0, 
/* out0042_em-eta2-phi23 */     0, 
/* out0043_em-eta0-phi22 */     1, 23, 3, 
/* out0044_em-eta0-phi23 */     0, 
/* out0045_em-eta15-phi-2 */     0, 
/* out0046_em-eta15-phi-1 */     0, 
/* out0047_em-eta15-phi0 */     1, 38, 1, 
/* out0048_em-eta15-phi1 */     0, 
/* out0049_em-eta16-phi-3 */     0, 
/* out0050_em-eta16-phi-1 */     1, 38, 1, 
/* out0051_em-eta16-phi0 */     1, 38, 1, 
/* out0052_em-eta16-phi2 */     0, 
/* out0053_em-eta16-phi4 */     0, 
/* out0054_em-eta16-phi5 */     0, 
/* out0055_em-eta16-phi6 */     0, 
/* out0056_em-eta16-phi7 */     0, 
/* out0057_em-eta17-phi5 */     0, 
/* out0058_em-eta17-phi6 */     0, 
/* out0059_em-eta17-phi7 */     0, 
/* out0060_em-eta17-phi8 */     0, 
/* out0061_em-eta15-phi10 */     1, 6, 1, 
/* out0062_em-eta15-phi11 */     1, 6, 1, 
/* out0063_em-eta15-phi12 */     1, 6, 1, 
/* out0064_em-eta15-phi13 */     1, 6, 1, 
/* out0065_em-eta16-phi10 */     1, 6, 1, 
/* out0066_em-eta16-phi12 */     1, 6, 1, 
/* out0067_em-eta16-phi13 */     1, 6, 1, 
/* out0068_em-eta17-phi12 */     0, 
/* out0069_em-eta12-phi14 */     1, 94, 1, 
/* out0070_em-eta12-phi15 */     1, 94, 1, 
/* out0071_em-eta12-phi16 */     0, 
/* out0072_em-eta13-phi14 */     1, 91, 1, 
/* out0073_em-eta13-phi15 */     1, 91, 1, 
/* out0074_em-eta13-phi16 */     1, 91, 1, 
/* out0075_em-eta13-phi17 */     0, 
/* out0076_em-eta14-phi16 */     1, 91, 1, 
/* out0077_em-eta9-phi17 */     1, 95, 1, 
/* out0078_em-eta9-phi18 */     1, 93, 1, 
/* out0079_em-eta10-phi16 */     1, 95, 1, 
/* out0080_em-eta10-phi17 */     1, 92, 1, 
/* out0081_em-eta10-phi18 */     1, 92, 1, 
/* out0082_em-eta10-phi19 */     1, 93, 1, 
/* out0083_em-eta11-phi17 */     1, 92, 1, 
/* out0084_em-eta11-phi18 */     1, 92, 1, 
/* out0085_em-eta7-phi18 */     4, 9, 1, 27, 2, 60, 2, 124, 2, 
/* out0086_em-eta7-phi19 */     0, 
/* out0087_em-eta8-phi18 */     2, 93, 1, 124, 1, 
/* out0088_em-eta8-phi19 */     1, 93, 2, 
/* out0089_em-eta8-phi20 */     3, 59, 1, 93, 1, 110, 1, 
/* out0090_em-eta9-phi19 */     1, 93, 1, 
/* out0091_em-eta5-phi19 */     4, 10, 1, 28, 2, 61, 2, 125, 2, 
/* out0092_em-eta5-phi20 */     0, 
/* out0093_em-eta6-phi19 */     1, 125, 1, 
/* out0094_em-eta6-phi20 */     0, 
/* out0095_em-eta3-phi20 */     5, 11, 1, 29, 2, 62, 1, 126, 1, 127, 2, 
/* out0096_em-eta4-phi20 */     2, 62, 1, 126, 1, 
/* out0097_em-eta2-phi20 */     6, 11, 1, 12, 2, 30, 3, 63, 4, 127, 3, 128, 1, 
/* out0098_em-eta2-phi21 */     1, 22, 2, 
/* out0099_em-eta0-phi21 */     2, 23, 5, 31, 1, 
/* out0100_em-eta1-phi21 */     4, 22, 5, 31, 1, 64, 1, 128, 1, 
/* out0101_em-eta11-phi-1 */     0, 
/* out0102_em-eta11-phi0 */     1, 39, 1, 
/* out0103_em-eta11-phi1 */     1, 117, 1, 
/* out0104_em-eta12-phi-2 */     1, 39, 1, 
/* out0105_em-eta12-phi-1 */     1, 39, 1, 
/* out0106_em-eta12-phi0 */     1, 39, 1, 
/* out0107_em-eta12-phi1 */     1, 39, 1, 
/* out0108_em-eta13-phi0 */     1, 39, 1, 
/* out0109_em-eta12-phi2 */     1, 117, 1, 
/* out0110_em-eta12-phi3 */     1, 117, 1, 
/* out0111_em-eta12-phi4 */     0, 
/* out0112_em-eta13-phi2 */     0, 
/* out0113_em-eta13-phi3 */     1, 116, 1, 
/* out0114_em-eta13-phi4 */     1, 116, 1, 
/* out0115_em-eta13-phi5 */     0, 
/* out0116_em-eta14-phi3 */     1, 116, 1, 
/* out0117_em-eta12-phi7 */     1, 7, 1, 
/* out0118_em-eta12-phi8 */     2, 7, 1, 65, 1, 
/* out0119_em-eta12-phi9 */     1, 65, 1, 
/* out0120_em-eta13-phi6 */     1, 7, 1, 
/* out0121_em-eta13-phi7 */     1, 7, 1, 
/* out0122_em-eta13-phi8 */     1, 7, 1, 
/* out0123_em-eta13-phi9 */     1, 7, 1, 
/* out0124_em-eta14-phi7 */     0, 
/* out0125_em-eta11-phi11 */     1, 8, 1, 
/* out0126_em-eta11-phi12 */     1, 8, 1, 
/* out0127_em-eta12-phi10 */     1, 8, 1, 
/* out0128_em-eta12-phi11 */     1, 8, 1, 
/* out0129_em-eta12-phi12 */     1, 8, 1, 
/* out0130_em-eta12-phi13 */     1, 8, 1, 
/* out0131_em-eta13-phi11 */     1, 8, 1, 
/* out0132_em-eta13-phi12 */     1, 8, 1, 
/* out0133_em-eta9-phi13 */     2, 14, 1, 97, 1, 
/* out0134_em-eta9-phi14 */     1, 97, 1, 
/* out0135_em-eta9-phi15 */     1, 95, 1, 
/* out0136_em-eta10-phi13 */     1, 94, 1, 
/* out0137_em-eta10-phi14 */     1, 94, 1, 
/* out0138_em-eta10-phi15 */     1, 94, 1, 
/* out0139_em-eta11-phi14 */     1, 94, 1, 
/* out0140_em-eta11-phi15 */     1, 94, 1, 
/* out0141_em-eta7-phi15 */     2, 98, 2, 111, 2, 
/* out0142_em-eta7-phi16 */     2, 98, 2, 111, 2, 
/* out0143_em-eta7-phi17 */     4, 9, 1, 27, 2, 60, 2, 124, 2, 
/* out0144_em-eta8-phi15 */     2, 95, 1, 97, 1, 
/* out0145_em-eta8-phi16 */     1, 95, 2, 
/* out0146_em-eta8-phi17 */     2, 95, 1, 124, 1, 
/* out0147_em-eta9-phi16 */     1, 95, 1, 
/* out0148_em-eta5-phi17 */     3, 9, 1, 41, 2, 66, 3, 
/* out0149_em-eta5-phi18 */     5, 9, 1, 10, 1, 28, 2, 61, 3, 125, 3, 
/* out0150_em-eta6-phi17 */     4, 9, 2, 27, 2, 60, 2, 124, 1, 
/* out0151_em-eta6-phi18 */     6, 9, 2, 27, 2, 60, 2, 61, 1, 124, 1, 125, 2, 
/* out0152_em-eta3-phi18 */     5, 11, 1, 45, 2, 46, 1, 129, 1, 130, 3, 
/* out0153_em-eta3-phi19 */     6, 11, 3, 29, 4, 62, 4, 126, 2, 127, 1, 130, 1, 
/* out0154_em-eta4-phi18 */     6, 10, 3, 28, 2, 45, 1, 61, 1, 126, 1, 129, 3, 
/* out0155_em-eta4-phi19 */     6, 10, 3, 28, 2, 29, 1, 61, 1, 62, 2, 126, 3, 
/* out0156_em-eta2-phi19 */     9, 11, 2, 12, 1, 29, 1, 30, 2, 46, 2, 63, 3, 127, 2, 130, 1, 131, 2, 
/* out0157_em-eta1-phi19 */     5, 12, 2, 30, 1, 47, 5, 131, 4, 132, 2, 
/* out0158_em-eta1-phi20 */     6, 12, 3, 30, 2, 31, 3, 63, 1, 64, 5, 128, 6, 
/* out0159_em-eta0-phi20 */     3, 31, 3, 64, 2, 132, 2, 
/* out0160_em-eta8-phi-1 */     5, 0, 1, 32, 1, 40, 1, 48, 1, 67, 1, 
/* out0161_em-eta8-phi0 */     5, 0, 2, 32, 1, 40, 1, 48, 1, 67, 1, 
/* out0162_em-eta9-phi-1 */     2, 0, 1, 40, 1, 
/* out0163_em-eta9-phi0 */     2, 0, 1, 40, 1, 
/* out0164_em-eta9-phi1 */     3, 0, 1, 40, 1, 118, 1, 
/* out0165_em-eta10-phi-1 */     2, 0, 1, 40, 1, 
/* out0166_em-eta10-phi0 */     2, 0, 1, 40, 1, 
/* out0167_em-eta9-phi2 */     1, 118, 1, 
/* out0168_em-eta9-phi3 */     2, 33, 1, 99, 1, 
/* out0169_em-eta10-phi1 */     1, 117, 1, 
/* out0170_em-eta10-phi2 */     1, 117, 1, 
/* out0171_em-eta10-phi3 */     1, 117, 1, 
/* out0172_em-eta11-phi2 */     1, 117, 1, 
/* out0173_em-eta11-phi3 */     1, 117, 1, 
/* out0174_em-eta9-phi5 */     2, 33, 1, 99, 1, 
/* out0175_em-eta9-phi6 */     1, 100, 1, 
/* out0176_em-eta10-phi4 */     1, 99, 1, 
/* out0177_em-eta10-phi5 */     1, 96, 1, 
/* out0178_em-eta10-phi6 */     1, 96, 1, 
/* out0179_em-eta10-phi7 */     1, 100, 1, 
/* out0180_em-eta11-phi5 */     1, 96, 1, 
/* out0181_em-eta11-phi6 */     1, 96, 1, 
/* out0182_em-eta9-phi8 */     2, 13, 1, 100, 1, 
/* out0183_em-eta9-phi9 */     2, 13, 1, 68, 1, 
/* out0184_em-eta9-phi10 */     3, 13, 1, 14, 1, 68, 1, 
/* out0185_em-eta10-phi8 */     2, 13, 1, 65, 1, 
/* out0186_em-eta10-phi9 */     2, 13, 1, 65, 1, 
/* out0187_em-eta10-phi10 */     2, 13, 1, 65, 1, 
/* out0188_em-eta11-phi8 */     2, 13, 1, 65, 1, 
/* out0189_em-eta11-phi9 */     2, 13, 1, 65, 1, 
/* out0190_em-eta8-phi11 */     2, 14, 1, 101, 1, 
/* out0191_em-eta8-phi12 */     2, 14, 1, 101, 1, 
/* out0192_em-eta9-phi11 */     1, 14, 1, 
/* out0193_em-eta9-phi12 */     1, 14, 1, 
/* out0194_em-eta10-phi11 */     1, 14, 1, 
/* out0195_em-eta10-phi12 */     1, 14, 1, 
/* out0196_em-eta6-phi13 */     0, 
/* out0197_em-eta6-phi14 */     0, 
/* out0198_em-eta7-phi13 */     1, 97, 1, 
/* out0199_em-eta7-phi14 */     2, 97, 1, 111, 1, 
/* out0200_em-eta8-phi13 */     1, 97, 1, 
/* out0201_em-eta8-phi14 */     1, 97, 2, 
/* out0202_em-eta5-phi15 */     2, 102, 3, 112, 3, 
/* out0203_em-eta5-phi16 */     2, 41, 2, 66, 2, 
/* out0204_em-eta6-phi15 */     2, 98, 2, 111, 2, 
/* out0205_em-eta6-phi16 */     3, 66, 1, 98, 2, 111, 1, 
/* out0206_em-eta3-phi16 */     2, 42, 4, 69, 4, 
/* out0207_em-eta3-phi17 */     3, 42, 1, 45, 3, 129, 1, 
/* out0208_em-eta4-phi16 */     4, 41, 2, 42, 1, 66, 1, 69, 2, 
/* out0209_em-eta4-phi17 */     4, 41, 2, 45, 2, 66, 1, 129, 3, 
/* out0210_em-eta2-phi17 */     0, 
/* out0211_em-eta2-phi18 */     3, 46, 5, 130, 3, 131, 1, 
/* out0212_em-eta1-phi18 */     2, 47, 2, 131, 1, 
/* out0213_em-eta0-phi18 */     0, 
/* out0214_em-eta0-phi19 */     2, 47, 1, 132, 4, 
/* out0215_em-eta5-phi-1 */     3, 34, 2, 49, 2, 70, 2, 
/* out0216_em-eta5-phi0 */     3, 34, 2, 49, 3, 70, 3, 
/* out0217_em-eta6-phi-1 */     4, 32, 1, 48, 1, 67, 1, 70, 1, 
/* out0218_em-eta6-phi0 */     5, 32, 1, 48, 1, 49, 1, 67, 1, 70, 1, 
/* out0219_em-eta7-phi-1 */     3, 32, 2, 48, 2, 67, 2, 
/* out0220_em-eta7-phi0 */     3, 32, 2, 48, 2, 67, 2, 
/* out0221_em-eta6-phi1 */     0, 
/* out0222_em-eta6-phi2 */     2, 50, 1, 71, 1, 
/* out0223_em-eta7-phi1 */     0, 
/* out0224_em-eta7-phi2 */     1, 118, 1, 
/* out0225_em-eta7-phi3 */     2, 50, 2, 71, 2, 
/* out0226_em-eta8-phi1 */     1, 118, 2, 
/* out0227_em-eta8-phi2 */     1, 118, 2, 
/* out0228_em-eta7-phi4 */     3, 33, 1, 50, 1, 71, 1, 
/* out0229_em-eta7-phi5 */     3, 72, 2, 119, 2, 133, 2, 
/* out0230_em-eta8-phi3 */     3, 33, 1, 99, 1, 118, 1, 
/* out0231_em-eta8-phi4 */     2, 33, 2, 99, 2, 
/* out0232_em-eta8-phi5 */     4, 33, 1, 99, 1, 119, 1, 133, 1, 
/* out0233_em-eta9-phi4 */     2, 33, 1, 99, 1, 
/* out0234_em-eta7-phi6 */     3, 72, 2, 119, 2, 133, 2, 
/* out0235_em-eta7-phi7 */     1, 73, 2, 
/* out0236_em-eta7-phi8 */     1, 73, 2, 
/* out0237_em-eta8-phi6 */     3, 100, 1, 119, 1, 133, 1, 
/* out0238_em-eta8-phi7 */     1, 100, 2, 
/* out0239_em-eta8-phi8 */     2, 68, 1, 100, 1, 
/* out0240_em-eta9-phi7 */     1, 100, 1, 
/* out0241_em-eta6-phi9 */     1, 2, 1, 
/* out0242_em-eta6-phi10 */     0, 
/* out0243_em-eta7-phi9 */     1, 68, 1, 
/* out0244_em-eta7-phi10 */     1, 68, 1, 
/* out0245_em-eta8-phi9 */     1, 68, 1, 
/* out0246_em-eta8-phi10 */     1, 68, 2, 
/* out0247_em-eta5-phi11 */     2, 25, 2, 103, 2, 
/* out0248_em-eta5-phi12 */     2, 25, 2, 103, 3, 
/* out0249_em-eta6-phi11 */     3, 24, 2, 101, 1, 103, 1, 
/* out0250_em-eta6-phi12 */     3, 24, 2, 101, 1, 103, 1, 
/* out0251_em-eta7-phi11 */     2, 24, 2, 101, 2, 
/* out0252_em-eta7-phi12 */     2, 24, 2, 101, 2, 
/* out0253_em-eta4-phi13 */     0, 
/* out0254_em-eta4-phi14 */     4, 102, 1, 104, 1, 112, 1, 113, 1, 
/* out0255_em-eta5-phi13 */     0, 
/* out0256_em-eta5-phi14 */     2, 102, 2, 112, 2, 
/* out0257_em-eta3-phi14 */     3, 20, 2, 104, 4, 113, 4, 
/* out0258_em-eta3-phi15 */     5, 20, 1, 42, 2, 69, 1, 104, 2, 113, 2, 
/* out0259_em-eta4-phi15 */     4, 69, 1, 102, 2, 112, 2, 113, 1, 
/* out0260_em-eta2-phi15 */     4, 20, 2, 43, 4, 74, 4, 106, 1, 
/* out0261_em-eta2-phi16 */     2, 43, 2, 74, 3, 
/* out0262_em-eta1-phi16 */     1, 43, 1, 
/* out0263_em-eta1-phi17 */     0, 
/* out0264_em-eta0-phi17 */     0, 
/* out0265_em-eta3-phi0 */     3, 35, 3, 51, 3, 75, 3, 
/* out0266_em-eta4-phi-1 */     5, 34, 2, 35, 1, 49, 1, 51, 1, 75, 1, 
/* out0267_em-eta4-phi0 */     6, 34, 2, 35, 1, 49, 1, 51, 1, 70, 1, 75, 1, 
/* out0268_em-eta4-phi1 */     0, 
/* out0269_em-eta4-phi2 */     4, 52, 2, 54, 1, 76, 1, 81, 1, 
/* out0270_em-eta5-phi1 */     0, 
/* out0271_em-eta5-phi2 */     2, 52, 1, 76, 2, 
/* out0272_em-eta5-phi3 */     2, 52, 2, 76, 3, 
/* out0273_em-eta5-phi4 */     0, 
/* out0274_em-eta6-phi3 */     2, 50, 2, 71, 2, 
/* out0275_em-eta6-phi4 */     2, 50, 2, 71, 2, 
/* out0276_em-eta5-phi5 */     0, 
/* out0277_em-eta5-phi6 */     3, 77, 3, 120, 3, 134, 3, 
/* out0278_em-eta6-phi5 */     3, 72, 2, 119, 1, 133, 1, 
/* out0279_em-eta6-phi6 */     5, 72, 2, 119, 1, 120, 1, 133, 1, 134, 2, 
/* out0280_em-eta5-phi7 */     4, 2, 1, 77, 2, 120, 2, 134, 2, 
/* out0281_em-eta5-phi8 */     2, 2, 2, 78, 3, 
/* out0282_em-eta6-phi7 */     5, 2, 2, 73, 2, 77, 1, 120, 1, 134, 1, 
/* out0283_em-eta6-phi8 */     2, 2, 2, 73, 2, 
/* out0284_em-eta4-phi9 */     3, 3, 2, 78, 1, 83, 1, 
/* out0285_em-eta4-phi10 */     0, 
/* out0286_em-eta5-phi9 */     1, 78, 2, 
/* out0287_em-eta5-phi10 */     0, 
/* out0288_em-eta3-phi12 */     2, 26, 3, 105, 2, 
/* out0289_em-eta4-phi11 */     2, 25, 2, 105, 2, 
/* out0290_em-eta4-phi12 */     3, 25, 2, 103, 1, 105, 2, 
/* out0291_em-eta2-phi13 */     2, 106, 1, 114, 1, 
/* out0292_em-eta3-phi13 */     0, 
/* out0293_em-eta2-phi14 */     5, 20, 3, 21, 1, 104, 1, 106, 4, 114, 5, 
/* out0294_em-eta1-phi15 */     5, 21, 1, 43, 1, 44, 4, 74, 1, 79, 5, 
/* out0295_em-eta0-phi16 */     0, 
/* out0296_em-eta2-phi-1 */     3, 36, 2, 53, 3, 80, 3, 
/* out0297_em-eta2-phi0 */     3, 36, 2, 53, 3, 80, 3, 
/* out0298_em-eta3-phi-1 */     3, 35, 3, 51, 3, 75, 3, 
/* out0299_em-eta2-phi1 */     2, 56, 1, 85, 1, 
/* out0300_em-eta3-phi1 */     0, 
/* out0301_em-eta3-phi2 */     2, 54, 4, 81, 4, 
/* out0302_em-eta3-phi3 */     2, 54, 2, 81, 2, 
/* out0303_em-eta4-phi3 */     2, 52, 3, 76, 2, 
/* out0304_em-eta3-phi4 */     0, 
/* out0305_em-eta3-phi5 */     1, 15, 3, 
/* out0306_em-eta4-phi4 */     0, 
/* out0307_em-eta4-phi5 */     0, 
/* out0308_em-eta3-phi6 */     1, 15, 3, 
/* out0309_em-eta3-phi7 */     5, 82, 4, 121, 2, 122, 1, 135, 2, 136, 1, 
/* out0310_em-eta4-phi6 */     3, 77, 1, 121, 1, 135, 1, 
/* out0311_em-eta4-phi7 */     5, 77, 1, 82, 2, 120, 1, 121, 3, 135, 3, 
/* out0312_em-eta3-phi8 */     8, 3, 2, 4, 1, 82, 1, 83, 2, 121, 1, 122, 1, 135, 1, 136, 2, 
/* out0313_em-eta3-phi9 */     3, 3, 1, 4, 1, 83, 4, 
/* out0314_em-eta4-phi8 */     5, 3, 3, 78, 2, 82, 1, 121, 1, 135, 1, 
/* out0315_em-eta2-phi10 */     1, 87, 1, 
/* out0316_em-eta3-phi10 */     0, 
/* out0317_em-eta3-phi11 */     2, 26, 3, 105, 2, 
/* out0318_em-eta2-phi11 */     2, 26, 1, 107, 3, 
/* out0319_em-eta2-phi12 */     2, 26, 1, 107, 3, 
/* out0320_em-eta1-phi12 */     3, 1, 1, 107, 1, 109, 3, 
/* out0321_em-eta1-phi13 */     4, 1, 2, 21, 1, 108, 1, 115, 2, 
/* out0322_em-eta0-phi14 */     2, 108, 3, 115, 2, 
/* out0323_em-eta1-phi14 */     7, 21, 5, 44, 1, 79, 1, 106, 2, 108, 3, 114, 2, 115, 3, 
/* out0324_em-eta0-phi15 */     2, 44, 3, 79, 2, 
/* out0325_em-eta1-phi-1 */     6, 36, 2, 37, 1, 53, 1, 55, 2, 80, 1, 84, 2, 
/* out0326_em-eta1-phi0 */     6, 36, 2, 37, 1, 53, 1, 55, 2, 80, 1, 84, 3, 
/* out0327_em-eta1-phi1 */     3, 56, 1, 57, 1, 88, 1, 
/* out0328_em-eta2-phi2 */     4, 54, 1, 56, 3, 81, 1, 85, 4, 
/* out0329_em-eta2-phi3 */     1, 16, 2, 
/* out0330_em-eta2-phi4 */     2, 16, 1, 17, 1, 
/* out0331_em-eta2-phi5 */     2, 15, 1, 17, 3, 
/* out0332_em-eta2-phi6 */     1, 15, 1, 
/* out0333_em-eta2-phi7 */     3, 86, 3, 122, 2, 136, 2, 
/* out0334_em-eta2-phi8 */     6, 4, 2, 86, 4, 122, 4, 123, 1, 136, 3, 137, 1, 
/* out0335_em-eta2-phi9 */     3, 4, 4, 83, 1, 87, 4, 
/* out0336_em-eta1-phi10 */     2, 5, 1, 90, 1, 
/* out0337_em-eta1-phi11 */     2, 107, 1, 109, 3, 
/* out0338_em-eta0-phi12 */     2, 1, 2, 109, 1, 
/* out0339_em-eta0-phi13 */     3, 1, 3, 108, 1, 115, 1, 
/* out0340_em-eta0-phi0 */     3, 37, 3, 55, 2, 84, 2, 
/* out0341_em-eta0-phi1 */     2, 57, 2, 88, 2, 
/* out0342_em-eta0-phi2 */     3, 18, 1, 57, 3, 88, 3, 
/* out0343_em-eta1-phi2 */     4, 56, 3, 57, 2, 85, 3, 88, 2, 
/* out0344_em-eta1-phi3 */     2, 16, 3, 18, 1, 
/* out0345_em-eta1-phi4 */     3, 16, 2, 17, 1, 19, 2, 
/* out0346_em-eta1-phi5 */     2, 17, 3, 19, 1, 
/* out0347_em-eta1-phi6 */     0, 
/* out0348_em-eta1-phi7 */     0, 
/* out0349_em-eta1-phi8 */     5, 5, 1, 86, 1, 89, 5, 123, 6, 137, 6, 
/* out0350_em-eta0-phi9 */     2, 5, 1, 90, 3, 
/* out0351_em-eta1-phi9 */     6, 5, 5, 87, 3, 89, 1, 90, 2, 123, 1, 137, 1, 
/* out0352_em-eta0-phi10 */     1, 90, 2, 
/* out0353_em-eta0-phi11 */     1, 109, 1, 
/* out0354_em-eta0-phi3 */     1, 18, 6, 
/* out0355_em-eta0-phi4 */     1, 19, 4, 
/* out0356_em-eta0-phi5 */     1, 19, 1, 
/* out0357_em-eta0-phi6 */     0, 
/* out0358_em-eta0-phi7 */     0, 
/* out0359_em-eta0-phi8 */     1, 89, 2, 
/* out0360_em-eta17-phi19 */     0, 
/* out0361_em-eta17-phi20 */     0, 
/* out0362_em-eta16-phi-2 */     1, 38, 1, 
/* out0363_em-eta16-phi1 */     1, 38, 1, 
/* out0364_em-eta17-phi0 */     1, 38, 1, 
/* out0365_em-eta17-phi3 */     0, 
/* out0366_em-eta17-phi4 */     0, 
/* out0367_em-eta16-phi11 */     1, 6, 1, 
/* out0368_em-eta14-phi14 */     1, 91, 1, 
/* out0369_em-eta14-phi15 */     1, 91, 1, 
/* out0370_em-eta11-phi16 */     1, 92, 1, 
/* out0371_em-eta13-phi-1 */     1, 39, 1, 
/* out0372_em-eta14-phi8 */     0, 
/* out0373_em-eta14-phi9 */     1, 7, 1, 
/* out0374_em-eta9-phi-2 */     1, 40, 1, 
/* out0375_em-eta11-phi7 */     1, 96, 1, 
/* out0376_em-eta14-phi19 */     0, 
/* out0377_em-eta14-phi17 */     1, 91, 1, 
/* out0378_em-eta11-phi19 */     1, 92, 1, 
/* out0379_em-eta14-phi4 */     1, 116, 1, 
/* out0380_em-eta14-phi6 */     1, 7, 1, 
/* out0381_em-eta11-phi4 */     1, 96, 1, 
/* out0382_em-eta14-phi21 */     0, 
/* out0383_em-eta11-phi22 */     1, 58, 1, 
/* out0384_em-eta12-phi17 */     1, 92, 1, 
/* out0385_em-eta14-phi2 */     1, 116, 1, 
/* out0386_em-eta11-phi13 */     1, 94, 1, 
/* out0387_em-eta12-phi6 */     1, 96, 1, 
/* out0388_em-eta11-phi10 */     1, 65, 1, 
/* out0389_em-eta4-phi23 */     0, 
/* out0390_em-eta17-phi11 */     0, 
/* out0391_em-eta12-phi18 */     1, 92, 1, 
/* out0392_em-eta12-phi5 */     1, 96, 1, 
/* out0393_em-eta0-phi-1 */     3, 37, 3, 55, 2, 84, 1, 
/* out0394_em-eta14-phi18 */     0, 
/* out0395_em-eta6-phi23 */     0, 
/* out0396_em-eta17-phi13 */     0, 
/* out0397_em-eta14-phi5 */     1, 116, 1, 
/* out0398_em-eta17-phi2 */     0, 
/* out0399_em-eta17-phi-2 */     1, 38, 1, 
/* out0400_em-eta17-phi1 */     1, 38, 1, 
/* out0401_em-eta17-phi10 */     0, 
/* out0402_em-eta15-phi15 */     0, 
/* out0403_em-eta14-phi0 */     1, 39, 1, 
/* out0404_em-eta15-phi8 */     0, 
/* out0405_em-eta13-phi10 */     0, 
/* out0406_em-eta13-phi13 */     0, 
/* out0407_em-eta15-phi20 */     0, 
/* out0408_em-eta17-phi-3 */     0, 
/* out0409_em-eta17-phi-1 */     0, 
/* out0410_em-eta15-phi16 */     1, 91, 1, 
/* out0411_em-eta13-phi-2 */     0, 
/* out0412_em-eta13-phi1 */     0, 
/* out0413_em-eta15-phi3 */     0, 
/* out0414_em-eta15-phi7 */     0, 
/* out0415_em-eta14-phi11 */     0, 
/* out0416_em-eta14-phi12 */     0, 
/* out0417_em-eta14-phi-1 */     0, 
/* out0418_em-eta15-phi14 */     0, 
/* out0419_em-eta15-phi9 */     0, 
/* out0420_em-eta10-phi-2 */     0, 
/* out0421_em-eta15-phi19 */     0, 
/* out0422_em-eta15-phi21 */     0, 
/* out0423_em-eta15-phi17 */     0, 
/* out0424_em-eta15-phi2 */     1, 116, 1, 
/* out0425_em-eta15-phi4 */     1, 116, 1, 
/* out0426_em-eta15-phi6 */     0, 
/* out0427_em-eta12-phi22 */     0
};