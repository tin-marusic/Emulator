parameter integer matrixE [0:1019] = {
/* num inputs = 63 (in0-in62) */
/* num outputs = 428 (out0-out427) */
/* max inputs per outputs = 5 */

/* out0_em-eta16-phi16 */     0, 
/* out1_em-eta16-phi17 */     1, 11, 1, 
/* out2_em-eta16-phi18 */     1, 11, 1, 
/* out3_em-eta16-phi19 */     0, 
/* out4_em-eta17-phi15 */     0, 
/* out5_em-eta17-phi16 */     1, 11, 1, 
/* out6_em-eta17-phi17 */     1, 11, 1, 
/* out7_em-eta17-phi18 */     1, 11, 1, 
/* out8_em-eta12-phi19 */     1, 9, 1, 
/* out9_em-eta12-phi20 */     1, 9, 1, 
/* out10_em-eta12-phi21 */     1, 9, 1, 
/* out11_em-eta13-phi18 */     1, 9, 1, 
/* out12_em-eta13-phi19 */     1, 9, 1, 
/* out13_em-eta13-phi20 */     1, 9, 1, 
/* out14_em-eta13-phi21 */     1, 9, 1, 
/* out15_em-eta14-phi20 */     1, 9, 1, 
/* out16_em-eta9-phi20 */     2, 10, 1, 25, 1, 
/* out17_em-eta9-phi21 */     1, 10, 1, 
/* out18_em-eta9-phi22 */     1, 10, 1, 
/* out19_em-eta10-phi20 */     1, 10, 1, 
/* out20_em-eta10-phi21 */     1, 10, 1, 
/* out21_em-eta10-phi22 */     1, 10, 1, 
/* out22_em-eta11-phi20 */     1, 10, 1, 
/* out23_em-eta11-phi21 */     1, 10, 1, 
/* out24_em-eta6-phi21 */     0, 
/* out25_em-eta6-phi22 */     0, 
/* out26_em-eta7-phi20 */     0, 
/* out27_em-eta7-phi21 */     0, 
/* out28_em-eta7-phi22 */     0, 
/* out29_em-eta8-phi21 */     0, 
/* out30_em-eta8-phi22 */     0, 
/* out31_em-eta4-phi21 */     0, 
/* out32_em-eta4-phi22 */     0, 
/* out33_em-eta5-phi21 */     0, 
/* out34_em-eta5-phi22 */     0, 
/* out35_em-eta5-phi23 */     0, 
/* out36_em-eta2-phi22 */     0, 
/* out37_em-eta3-phi21 */     0, 
/* out38_em-eta3-phi22 */     0, 
/* out39_em-eta3-phi23 */     0, 
/* out40_em-eta1-phi22 */     0, 
/* out41_em-eta1-phi23 */     0, 
/* out42_em-eta2-phi23 */     0, 
/* out43_em-eta0-phi22 */     0, 
/* out44_em-eta0-phi23 */     0, 
/* out45_em-eta15-phi-2 */     0, 
/* out46_em-eta15-phi-1 */     0, 
/* out47_em-eta15-phi0 */     0, 
/* out48_em-eta15-phi1 */     0, 
/* out49_em-eta16-phi-3 */     0, 
/* out50_em-eta16-phi-1 */     0, 
/* out51_em-eta16-phi0 */     0, 
/* out52_em-eta16-phi2 */     0, 
/* out53_em-eta16-phi4 */     0, 
/* out54_em-eta16-phi5 */     1, 19, 1, 
/* out55_em-eta16-phi6 */     1, 19, 1, 
/* out56_em-eta16-phi7 */     0, 
/* out57_em-eta17-phi5 */     1, 19, 1, 
/* out58_em-eta17-phi6 */     1, 19, 1, 
/* out59_em-eta17-phi7 */     1, 19, 1, 
/* out60_em-eta17-phi8 */     0, 
/* out61_em-eta15-phi10 */     0, 
/* out62_em-eta15-phi11 */     0, 
/* out63_em-eta15-phi12 */     0, 
/* out64_em-eta15-phi13 */     0, 
/* out65_em-eta16-phi10 */     0, 
/* out66_em-eta16-phi12 */     0, 
/* out67_em-eta16-phi13 */     0, 
/* out68_em-eta17-phi12 */     0, 
/* out69_em-eta12-phi14 */     0, 
/* out70_em-eta12-phi15 */     0, 
/* out71_em-eta12-phi16 */     0, 
/* out72_em-eta13-phi14 */     0, 
/* out73_em-eta13-phi15 */     0, 
/* out74_em-eta13-phi16 */     0, 
/* out75_em-eta13-phi17 */     0, 
/* out76_em-eta14-phi16 */     0, 
/* out77_em-eta9-phi17 */     1, 26, 1, 
/* out78_em-eta9-phi18 */     1, 25, 1, 
/* out79_em-eta10-phi16 */     0, 
/* out80_em-eta10-phi17 */     1, 24, 1, 
/* out81_em-eta10-phi18 */     1, 24, 1, 
/* out82_em-eta10-phi19 */     0, 
/* out83_em-eta11-phi17 */     1, 24, 1, 
/* out84_em-eta11-phi18 */     1, 24, 1, 
/* out85_em-eta7-phi18 */     2, 13, 1, 49, 2, 
/* out86_em-eta7-phi19 */     1, 25, 1, 
/* out87_em-eta8-phi18 */     2, 25, 1, 49, 1, 
/* out88_em-eta8-phi19 */     1, 25, 2, 
/* out89_em-eta8-phi20 */     1, 25, 1, 
/* out90_em-eta9-phi19 */     1, 25, 1, 
/* out91_em-eta5-phi19 */     2, 14, 1, 50, 2, 
/* out92_em-eta5-phi20 */     0, 
/* out93_em-eta6-phi19 */     1, 50, 1, 
/* out94_em-eta6-phi20 */     0, 
/* out95_em-eta3-phi20 */     3, 15, 1, 51, 1, 52, 2, 
/* out96_em-eta4-phi20 */     1, 51, 1, 
/* out97_em-eta2-phi20 */     4, 15, 1, 16, 2, 52, 3, 53, 1, 
/* out98_em-eta2-phi21 */     0, 
/* out99_em-eta0-phi21 */     0, 
/* out100_em-eta1-phi21 */     1, 53, 1, 
/* out101_em-eta11-phi-1 */     0, 
/* out102_em-eta11-phi0 */     0, 
/* out103_em-eta11-phi1 */     0, 
/* out104_em-eta12-phi-2 */     0, 
/* out105_em-eta12-phi-1 */     0, 
/* out106_em-eta12-phi0 */     0, 
/* out107_em-eta12-phi1 */     0, 
/* out108_em-eta13-phi0 */     0, 
/* out109_em-eta12-phi2 */     0, 
/* out110_em-eta12-phi3 */     1, 12, 1, 
/* out111_em-eta12-phi4 */     1, 12, 1, 
/* out112_em-eta13-phi2 */     1, 12, 1, 
/* out113_em-eta13-phi3 */     1, 12, 1, 
/* out114_em-eta13-phi4 */     1, 12, 1, 
/* out115_em-eta13-phi5 */     1, 12, 1, 
/* out116_em-eta14-phi3 */     1, 12, 1, 
/* out117_em-eta12-phi7 */     0, 
/* out118_em-eta12-phi8 */     0, 
/* out119_em-eta12-phi9 */     0, 
/* out120_em-eta13-phi6 */     0, 
/* out121_em-eta13-phi7 */     0, 
/* out122_em-eta13-phi8 */     0, 
/* out123_em-eta13-phi9 */     0, 
/* out124_em-eta14-phi7 */     0, 
/* out125_em-eta11-phi11 */     0, 
/* out126_em-eta11-phi12 */     0, 
/* out127_em-eta12-phi10 */     0, 
/* out128_em-eta12-phi11 */     0, 
/* out129_em-eta12-phi12 */     0, 
/* out130_em-eta12-phi13 */     0, 
/* out131_em-eta13-phi11 */     0, 
/* out132_em-eta13-phi12 */     0, 
/* out133_em-eta9-phi13 */     0, 
/* out134_em-eta9-phi14 */     0, 
/* out135_em-eta9-phi15 */     1, 26, 1, 
/* out136_em-eta10-phi13 */     0, 
/* out137_em-eta10-phi14 */     0, 
/* out138_em-eta10-phi15 */     0, 
/* out139_em-eta11-phi14 */     0, 
/* out140_em-eta11-phi15 */     0, 
/* out141_em-eta7-phi15 */     0, 
/* out142_em-eta7-phi16 */     1, 26, 1, 
/* out143_em-eta7-phi17 */     2, 13, 1, 49, 2, 
/* out144_em-eta8-phi15 */     1, 26, 1, 
/* out145_em-eta8-phi16 */     1, 26, 2, 
/* out146_em-eta8-phi17 */     2, 26, 1, 49, 1, 
/* out147_em-eta9-phi16 */     1, 26, 1, 
/* out148_em-eta5-phi17 */     1, 13, 1, 
/* out149_em-eta5-phi18 */     3, 13, 1, 14, 1, 50, 3, 
/* out150_em-eta6-phi17 */     2, 13, 2, 49, 1, 
/* out151_em-eta6-phi18 */     3, 13, 2, 49, 1, 50, 2, 
/* out152_em-eta3-phi18 */     2, 0, 2, 15, 1, 
/* out153_em-eta3-phi19 */     3, 15, 3, 51, 2, 52, 1, 
/* out154_em-eta4-phi18 */     2, 14, 3, 51, 1, 
/* out155_em-eta4-phi19 */     2, 14, 3, 51, 3, 
/* out156_em-eta2-phi19 */     4, 1, 1, 15, 2, 16, 1, 52, 2, 
/* out157_em-eta1-phi19 */     3, 1, 1, 2, 1, 16, 2, 
/* out158_em-eta1-phi20 */     2, 16, 3, 53, 6, 
/* out159_em-eta0-phi20 */     0, 
/* out160_em-eta8-phi-1 */     0, 
/* out161_em-eta8-phi0 */     0, 
/* out162_em-eta9-phi-1 */     0, 
/* out163_em-eta9-phi0 */     0, 
/* out164_em-eta9-phi1 */     1, 17, 1, 
/* out165_em-eta10-phi-1 */     0, 
/* out166_em-eta10-phi0 */     0, 
/* out167_em-eta9-phi2 */     1, 17, 1, 
/* out168_em-eta9-phi3 */     1, 17, 1, 
/* out169_em-eta10-phi1 */     1, 17, 1, 
/* out170_em-eta10-phi2 */     1, 17, 1, 
/* out171_em-eta10-phi3 */     1, 17, 1, 
/* out172_em-eta11-phi2 */     1, 17, 1, 
/* out173_em-eta11-phi3 */     1, 17, 1, 
/* out174_em-eta9-phi5 */     0, 
/* out175_em-eta9-phi6 */     0, 
/* out176_em-eta10-phi4 */     0, 
/* out177_em-eta10-phi5 */     0, 
/* out178_em-eta10-phi6 */     0, 
/* out179_em-eta10-phi7 */     0, 
/* out180_em-eta11-phi5 */     0, 
/* out181_em-eta11-phi6 */     0, 
/* out182_em-eta9-phi8 */     0, 
/* out183_em-eta9-phi9 */     0, 
/* out184_em-eta9-phi10 */     0, 
/* out185_em-eta10-phi8 */     0, 
/* out186_em-eta10-phi9 */     0, 
/* out187_em-eta10-phi10 */     0, 
/* out188_em-eta11-phi8 */     0, 
/* out189_em-eta11-phi9 */     0, 
/* out190_em-eta8-phi11 */     1, 54, 2, 
/* out191_em-eta8-phi12 */     1, 54, 2, 
/* out192_em-eta9-phi11 */     0, 
/* out193_em-eta9-phi12 */     0, 
/* out194_em-eta10-phi11 */     0, 
/* out195_em-eta10-phi12 */     0, 
/* out196_em-eta6-phi13 */     1, 20, 2, 
/* out197_em-eta6-phi14 */     1, 20, 1, 
/* out198_em-eta7-phi13 */     0, 
/* out199_em-eta7-phi14 */     0, 
/* out200_em-eta8-phi13 */     0, 
/* out201_em-eta8-phi14 */     0, 
/* out202_em-eta5-phi15 */     0, 
/* out203_em-eta5-phi16 */     0, 
/* out204_em-eta6-phi15 */     0, 
/* out205_em-eta6-phi16 */     0, 
/* out206_em-eta3-phi16 */     0, 
/* out207_em-eta3-phi17 */     1, 0, 2, 
/* out208_em-eta4-phi16 */     0, 
/* out209_em-eta4-phi17 */     0, 
/* out210_em-eta2-phi17 */     2, 0, 2, 3, 2, 
/* out211_em-eta2-phi18 */     2, 0, 2, 1, 2, 
/* out212_em-eta1-phi18 */     2, 1, 4, 4, 1, 
/* out213_em-eta0-phi18 */     2, 2, 2, 4, 3, 
/* out214_em-eta0-phi19 */     1, 2, 5, 
/* out215_em-eta5-phi-1 */     0, 
/* out216_em-eta5-phi0 */     0, 
/* out217_em-eta6-phi-1 */     0, 
/* out218_em-eta6-phi0 */     2, 27, 1, 40, 1, 
/* out219_em-eta7-phi-1 */     0, 
/* out220_em-eta7-phi0 */     0, 
/* out221_em-eta6-phi1 */     2, 27, 2, 40, 2, 
/* out222_em-eta6-phi2 */     3, 18, 1, 27, 1, 40, 2, 
/* out223_em-eta7-phi1 */     2, 18, 2, 40, 1, 
/* out224_em-eta7-phi2 */     1, 18, 2, 
/* out225_em-eta7-phi3 */     1, 18, 1, 
/* out226_em-eta8-phi1 */     1, 18, 1, 
/* out227_em-eta8-phi2 */     1, 18, 1, 
/* out228_em-eta7-phi4 */     0, 
/* out229_em-eta7-phi5 */     0, 
/* out230_em-eta8-phi3 */     0, 
/* out231_em-eta8-phi4 */     0, 
/* out232_em-eta8-phi5 */     0, 
/* out233_em-eta9-phi4 */     0, 
/* out234_em-eta7-phi6 */     0, 
/* out235_em-eta7-phi7 */     1, 35, 1, 
/* out236_em-eta7-phi8 */     1, 35, 1, 
/* out237_em-eta8-phi6 */     0, 
/* out238_em-eta8-phi7 */     0, 
/* out239_em-eta8-phi8 */     0, 
/* out240_em-eta9-phi7 */     0, 
/* out241_em-eta6-phi9 */     2, 35, 1, 45, 2, 
/* out242_em-eta6-phi10 */     1, 45, 2, 
/* out243_em-eta7-phi9 */     1, 45, 1, 
/* out244_em-eta7-phi10 */     1, 45, 1, 
/* out245_em-eta8-phi9 */     0, 
/* out246_em-eta8-phi10 */     0, 
/* out247_em-eta5-phi11 */     1, 55, 2, 
/* out248_em-eta5-phi12 */     1, 55, 2, 
/* out249_em-eta6-phi11 */     2, 45, 1, 55, 2, 
/* out250_em-eta6-phi12 */     1, 55, 2, 
/* out251_em-eta7-phi11 */     1, 54, 2, 
/* out252_em-eta7-phi12 */     1, 54, 2, 
/* out253_em-eta4-phi13 */     1, 21, 3, 
/* out254_em-eta4-phi14 */     1, 21, 1, 
/* out255_em-eta5-phi13 */     1, 20, 3, 
/* out256_em-eta5-phi14 */     1, 20, 2, 
/* out257_em-eta3-phi14 */     0, 
/* out258_em-eta3-phi15 */     0, 
/* out259_em-eta4-phi15 */     0, 
/* out260_em-eta2-phi15 */     0, 
/* out261_em-eta2-phi16 */     1, 3, 1, 
/* out262_em-eta1-phi16 */     2, 3, 1, 5, 1, 
/* out263_em-eta1-phi17 */     2, 3, 4, 4, 1, 
/* out264_em-eta0-phi17 */     2, 4, 3, 5, 2, 
/* out265_em-eta3-phi0 */     1, 42, 1, 
/* out266_em-eta4-phi-1 */     0, 
/* out267_em-eta4-phi0 */     2, 28, 1, 41, 1, 
/* out268_em-eta4-phi1 */     2, 28, 3, 41, 3, 
/* out269_em-eta4-phi2 */     2, 28, 1, 41, 1, 
/* out270_em-eta5-phi1 */     3, 27, 2, 40, 1, 41, 2, 
/* out271_em-eta5-phi2 */     2, 27, 2, 40, 1, 
/* out272_em-eta5-phi3 */     0, 
/* out273_em-eta5-phi4 */     2, 29, 2, 56, 2, 
/* out274_em-eta6-phi3 */     0, 
/* out275_em-eta6-phi4 */     1, 56, 1, 
/* out276_em-eta5-phi5 */     2, 29, 2, 56, 3, 
/* out277_em-eta5-phi6 */     0, 
/* out278_em-eta6-phi5 */     1, 56, 2, 
/* out279_em-eta6-phi6 */     0, 
/* out280_em-eta5-phi7 */     0, 
/* out281_em-eta5-phi8 */     2, 35, 1, 36, 2, 
/* out282_em-eta6-phi7 */     1, 35, 2, 
/* out283_em-eta6-phi8 */     1, 35, 2, 
/* out284_em-eta4-phi9 */     2, 36, 2, 46, 1, 
/* out285_em-eta4-phi10 */     2, 6, 2, 46, 3, 
/* out286_em-eta5-phi9 */     1, 36, 1, 
/* out287_em-eta5-phi10 */     2, 45, 1, 46, 2, 
/* out288_em-eta3-phi12 */     2, 57, 1, 59, 1, 
/* out289_em-eta4-phi11 */     2, 46, 1, 57, 3, 
/* out290_em-eta4-phi12 */     2, 21, 1, 57, 3, 
/* out291_em-eta2-phi13 */     1, 22, 4, 
/* out292_em-eta3-phi13 */     2, 21, 3, 22, 1, 
/* out293_em-eta2-phi14 */     0, 
/* out294_em-eta1-phi15 */     0, 
/* out295_em-eta0-phi16 */     1, 5, 5, 
/* out296_em-eta2-phi-1 */     0, 
/* out297_em-eta2-phi0 */     3, 30, 2, 42, 1, 43, 1, 
/* out298_em-eta3-phi-1 */     0, 
/* out299_em-eta2-phi1 */     3, 30, 4, 42, 3, 43, 1, 
/* out300_em-eta3-phi1 */     4, 28, 2, 30, 1, 41, 1, 42, 3, 
/* out301_em-eta3-phi2 */     1, 28, 1, 
/* out302_em-eta3-phi3 */     3, 31, 2, 58, 1, 60, 2, 
/* out303_em-eta4-phi3 */     1, 58, 1, 
/* out304_em-eta3-phi4 */     3, 31, 4, 58, 2, 60, 1, 
/* out305_em-eta3-phi5 */     0, 
/* out306_em-eta4-phi4 */     3, 29, 2, 31, 1, 58, 3, 
/* out307_em-eta4-phi5 */     2, 29, 2, 58, 1, 
/* out308_em-eta3-phi6 */     0, 
/* out309_em-eta3-phi7 */     0, 
/* out310_em-eta4-phi6 */     0, 
/* out311_em-eta4-phi7 */     0, 
/* out312_em-eta3-phi8 */     1, 37, 2, 
/* out313_em-eta3-phi9 */     2, 6, 1, 37, 3, 
/* out314_em-eta4-phi8 */     1, 36, 3, 
/* out315_em-eta2-phi10 */     4, 6, 1, 7, 3, 47, 2, 48, 2, 
/* out316_em-eta3-phi10 */     3, 6, 3, 46, 1, 47, 4, 
/* out317_em-eta3-phi11 */     4, 6, 1, 47, 1, 57, 1, 59, 1, 
/* out318_em-eta2-phi11 */     4, 7, 2, 47, 1, 48, 1, 59, 3, 
/* out319_em-eta2-phi12 */     2, 22, 2, 59, 3, 
/* out320_em-eta1-phi12 */     1, 61, 4, 
/* out321_em-eta1-phi13 */     1, 22, 1, 
/* out322_em-eta0-phi14 */     0, 
/* out323_em-eta1-phi14 */     0, 
/* out324_em-eta0-phi15 */     0, 
/* out325_em-eta1-phi-1 */     0, 
/* out326_em-eta1-phi0 */     3, 23, 2, 32, 2, 43, 2, 
/* out327_em-eta1-phi1 */     4, 23, 3, 32, 4, 43, 4, 44, 1, 
/* out328_em-eta2-phi2 */     1, 30, 1, 
/* out329_em-eta2-phi3 */     3, 33, 3, 60, 3, 62, 1, 
/* out330_em-eta2-phi4 */     3, 31, 1, 33, 2, 60, 2, 
/* out331_em-eta2-phi5 */     0, 
/* out332_em-eta2-phi6 */     0, 
/* out333_em-eta2-phi7 */     0, 
/* out334_em-eta2-phi8 */     1, 37, 1, 
/* out335_em-eta2-phi9 */     2, 37, 2, 38, 3, 
/* out336_em-eta1-phi10 */     5, 7, 2, 8, 2, 38, 1, 39, 1, 48, 3, 
/* out337_em-eta1-phi11 */     4, 7, 1, 8, 1, 48, 2, 61, 3, 
/* out338_em-eta0-phi12 */     1, 61, 1, 
/* out339_em-eta0-phi13 */     0, 
/* out340_em-eta0-phi0 */     3, 23, 1, 32, 1, 44, 3, 
/* out341_em-eta0-phi1 */     3, 23, 2, 32, 1, 44, 4, 
/* out342_em-eta0-phi2 */     1, 34, 1, 
/* out343_em-eta1-phi2 */     1, 62, 1, 
/* out344_em-eta1-phi3 */     3, 33, 2, 34, 3, 62, 6, 
/* out345_em-eta1-phi4 */     1, 33, 1, 
/* out346_em-eta1-phi5 */     0, 
/* out347_em-eta1-phi6 */     0, 
/* out348_em-eta1-phi7 */     0, 
/* out349_em-eta1-phi8 */     0, 
/* out350_em-eta0-phi9 */     1, 39, 4, 
/* out351_em-eta1-phi9 */     2, 38, 4, 39, 1, 
/* out352_em-eta0-phi10 */     2, 8, 3, 39, 2, 
/* out353_em-eta0-phi11 */     1, 8, 2, 
/* out354_em-eta0-phi3 */     1, 34, 4, 
/* out355_em-eta0-phi4 */     0, 
/* out356_em-eta0-phi5 */     0, 
/* out357_em-eta0-phi6 */     0, 
/* out358_em-eta0-phi7 */     0, 
/* out359_em-eta0-phi8 */     0, 
/* out360_em-eta17-phi19 */     1, 11, 1, 
/* out361_em-eta17-phi20 */     1, 11, 1, 
/* out362_em-eta16-phi-2 */     0, 
/* out363_em-eta16-phi1 */     0, 
/* out364_em-eta17-phi0 */     0, 
/* out365_em-eta17-phi3 */     1, 19, 1, 
/* out366_em-eta17-phi4 */     1, 19, 1, 
/* out367_em-eta16-phi11 */     0, 
/* out368_em-eta14-phi14 */     0, 
/* out369_em-eta14-phi15 */     0, 
/* out370_em-eta11-phi16 */     1, 24, 1, 
/* out371_em-eta13-phi-1 */     0, 
/* out372_em-eta14-phi8 */     0, 
/* out373_em-eta14-phi9 */     0, 
/* out374_em-eta9-phi-2 */     0, 
/* out375_em-eta11-phi7 */     0, 
/* out376_em-eta14-phi19 */     0, 
/* out377_em-eta14-phi17 */     0, 
/* out378_em-eta11-phi19 */     1, 24, 1, 
/* out379_em-eta14-phi4 */     1, 12, 1, 
/* out380_em-eta14-phi6 */     0, 
/* out381_em-eta11-phi4 */     0, 
/* out382_em-eta14-phi21 */     0, 
/* out383_em-eta11-phi22 */     0, 
/* out384_em-eta12-phi17 */     1, 24, 1, 
/* out385_em-eta14-phi2 */     0, 
/* out386_em-eta11-phi13 */     0, 
/* out387_em-eta12-phi6 */     0, 
/* out388_em-eta11-phi10 */     0, 
/* out389_em-eta4-phi23 */     0, 
/* out390_em-eta17-phi11 */     0, 
/* out391_em-eta12-phi18 */     1, 24, 1, 
/* out392_em-eta12-phi5 */     0, 
/* out393_em-eta0-phi-1 */     0, 
/* out394_em-eta14-phi18 */     0, 
/* out395_em-eta6-phi23 */     0, 
/* out396_em-eta17-phi13 */     0, 
/* out397_em-eta14-phi5 */     0, 
/* out398_em-eta17-phi2 */     0, 
/* out399_em-eta17-phi-2 */     0, 
/* out400_em-eta17-phi1 */     0, 
/* out401_em-eta17-phi10 */     0, 
/* out402_em-eta15-phi15 */     0, 
/* out403_em-eta14-phi0 */     0, 
/* out404_em-eta15-phi8 */     0, 
/* out405_em-eta13-phi10 */     0, 
/* out406_em-eta13-phi13 */     0, 
/* out407_em-eta15-phi20 */     0, 
/* out408_em-eta17-phi-3 */     0, 
/* out409_em-eta17-phi-1 */     0, 
/* out410_em-eta15-phi16 */     0, 
/* out411_em-eta13-phi-2 */     0, 
/* out412_em-eta13-phi1 */     0, 
/* out413_em-eta15-phi3 */     0, 
/* out414_em-eta15-phi7 */     0, 
/* out415_em-eta14-phi11 */     0, 
/* out416_em-eta14-phi12 */     0, 
/* out417_em-eta14-phi-1 */     0, 
/* out418_em-eta15-phi14 */     0, 
/* out419_em-eta15-phi9 */     0, 
/* out420_em-eta10-phi-2 */     0, 
/* out421_em-eta15-phi19 */     0, 
/* out422_em-eta15-phi21 */     0, 
/* out423_em-eta15-phi17 */     0, 
/* out424_em-eta15-phi2 */     0, 
/* out425_em-eta15-phi4 */     0, 
/* out426_em-eta15-phi6 */     0, 
/* out427_em-eta12-phi22 */     0

};
