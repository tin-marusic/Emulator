parameter integer matrixH [0:2180] = {
/* num inputs = 157 (in0-in156) */
/* num outputs = 515(out0-out514) */
//* max inputs per outputs = 9 */
//* total number of input in adders 833 */

/* out0000_had-eta14-phi21 */     1, 118, 2, 
/* out0001_had-eta14-phi22 */     3, 78, 2, 107, 2, 118, 2, 
/* out0002_had-eta14-phi23 */     3, 78, 2, 107, 2, 118, 2, 
/* out0003_had-eta15-phi21 */     1, 77, 2, 
/* out0004_had-eta15-phi22 */     3, 77, 2, 107, 2, 118, 2, 
/* out0005_had-eta15-phi23 */     3, 77, 2, 107, 2, 118, 2, 
/* out0006_had-eta15-phi24 */     0, 
/* out0007_had-eta16-phi22 */     1, 77, 2, 
/* out0008_had-eta11-phi22 */     2, 108, 2, 119, 2, 
/* out0009_had-eta11-phi23 */     3, 79, 2, 108, 4, 119, 4, 
/* out0010_had-eta11-phi24 */     2, 108, 2, 119, 2, 
/* out0011_had-eta12-phi22 */     2, 78, 2, 119, 2, 
/* out0012_had-eta12-phi23 */     3, 78, 2, 108, 2, 119, 2, 
/* out0013_had-eta12-phi24 */     1, 78, 2, 
/* out0014_had-eta13-phi22 */     3, 78, 2, 107, 2, 118, 2, 
/* out0015_had-eta13-phi23 */     3, 78, 2, 107, 2, 118, 2, 
/* out0016_had-eta8-phi22 */     5, 96, 2, 109, 2, 120, 2, 137, 2, 139, 1, 
/* out0017_had-eta8-phi23 */     5, 109, 4, 120, 4, 121, 4, 137, 2, 139, 1, 
/* out0018_had-eta9-phi22 */     4, 79, 2, 96, 2, 109, 2, 120, 2, 
/* out0019_had-eta9-phi23 */     3, 79, 4, 109, 4, 120, 4, 
/* out0020_had-eta9-phi24 */     2, 109, 2, 120, 2, 
/* out0021_had-eta10-phi22 */     3, 79, 2, 108, 2, 119, 2, 
/* out0022_had-eta10-phi23 */     4, 79, 4, 108, 4, 119, 2, 120, 2, 
/* out0023_had-eta6-phi22 */     5, 80, 4, 100, 2, 110, 2, 137, 3, 139, 2, 
/* out0024_had-eta6-phi23 */     6, 80, 4, 110, 4, 111, 2, 121, 2, 137, 3, 139, 2, 
/* out0025_had-eta6-phi24 */     0, 
/* out0026_had-eta7-phi22 */     5, 80, 4, 110, 2, 121, 2, 137, 2, 139, 2, 
/* out0027_had-eta7-phi23 */     5, 80, 4, 110, 6, 121, 6, 137, 2, 139, 2, 
/* out0028_had-eta7-phi24 */     2, 110, 2, 121, 2, 
/* out0029_had-eta4-phi22 */     6, 81, 2, 82, 2, 101, 2, 102, 2, 138, 1, 140, 1, 
/* out0030_had-eta4-phi23 */     5, 81, 2, 82, 4, 111, 2, 138, 1, 140, 1, 
/* out0031_had-eta5-phi22 */     5, 81, 6, 101, 4, 111, 2, 137, 1, 139, 3, 
/* out0032_had-eta5-phi23 */     4, 81, 6, 111, 8, 137, 1, 139, 3, 
/* out0033_had-eta5-phi24 */     1, 111, 2, 
/* out0034_had-eta3-phi22 */     4, 82, 4, 102, 6, 138, 1, 140, 1, 
/* out0035_had-eta3-phi23 */     4, 82, 6, 83, 2, 138, 1, 140, 1, 
/* out0036_had-eta3-phi24 */     0, 
/* out0037_had-eta1-phi23 */     3, 84, 12, 138, 2, 140, 1, 
/* out0038_had-eta2-phi23 */     4, 83, 10, 84, 2, 138, 2, 140, 1, 
/* out0039_had-eta2-phi24 */     0, 
/* out0040_had-eta15-phi16 */     1, 112, 2, 
/* out0041_had-eta15-phi17 */     2, 30, 2, 112, 2, 
/* out0042_had-eta15-phi18 */     0, 
/* out0043_had-eta15-phi19 */     2, 30, 2, 94, 2, 
/* out0044_had-eta16-phi16 */     0, 
/* out0045_had-eta16-phi17 */     0, 
/* out0046_had-eta16-phi18 */     0, 
/* out0047_had-eta16-phi19 */     0, 
/* out0048_had-eta11-phi19 */     2, 31, 2, 95, 2, 
/* out0049_had-eta12-phi18 */     2, 31, 2, 125, 2, 
/* out0050_had-eta12-phi19 */     1, 31, 2, 
/* out0051_had-eta12-phi20 */     2, 31, 2, 95, 2, 
/* out0052_had-eta13-phi18 */     2, 30, 2, 94, 2, 
/* out0053_had-eta13-phi19 */     1, 94, 2, 
/* out0054_had-eta13-phi20 */     1, 94, 2, 
/* out0055_had-eta14-phi19 */     2, 30, 2, 94, 2, 
/* out0056_had-eta9-phi19 */     0, 
/* out0057_had-eta9-phi20 */     2, 96, 2, 99, 2, 
/* out0058_had-eta9-phi21 */     2, 96, 4, 99, 2, 
/* out0059_had-eta10-phi19 */     2, 31, 2, 95, 2, 
/* out0060_had-eta10-phi20 */     2, 31, 2, 95, 2, 
/* out0061_had-eta10-phi21 */     1, 95, 2, 
/* out0062_had-eta11-phi20 */     2, 31, 2, 95, 2, 
/* out0063_had-eta7-phi20 */     1, 99, 2, 
/* out0064_had-eta7-phi21 */     2, 99, 2, 100, 4, 
/* out0065_had-eta8-phi20 */     2, 96, 2, 99, 4, 
/* out0066_had-eta8-phi21 */     2, 96, 4, 99, 4, 
/* out0067_had-eta5-phi21 */     2, 100, 2, 101, 6, 
/* out0068_had-eta6-phi21 */     1, 100, 6, 
/* out0069_had-eta3-phi21 */     2, 102, 6, 131, 2, 
/* out0070_had-eta4-phi21 */     3, 101, 4, 102, 2, 131, 6, 
/* out0071_had-eta2-phi21 */     1, 132, 1, 
/* out0072_had-eta2-phi22 */     3, 83, 4, 138, 2, 140, 1, 
/* out0073_had-eta1-phi22 */     3, 84, 2, 138, 2, 140, 1, 
/* out0074_had-eta16-phi1 */     0, 
/* out0075_had-eta16-phi2 */     0, 
/* out0076_had-eta16-phi3 */     0, 
/* out0077_had-eta16-phi4 */     0, 
/* out0078_had-eta17-phi1 */     0, 
/* out0079_had-eta17-phi2 */     0, 
/* out0080_had-eta17-phi3 */     0, 
/* out0081_had-eta17-phi4 */     0, 
/* out0082_had-eta16-phi7 */     0, 
/* out0083_had-eta16-phi8 */     0, 
/* out0084_had-eta16-phi9 */     0, 
/* out0085_had-eta16-phi10 */     0, 
/* out0086_had-eta17-phi6 */     0, 
/* out0087_had-eta17-phi8 */     0, 
/* out0088_had-eta17-phi9 */     0, 
/* out0089_had-eta17-phi10 */     0, 
/* out0090_had-eta14-phi12 */     0, 
/* out0091_had-eta14-phi13 */     1, 32, 2, 
/* out0092_had-eta14-phi14 */     1, 32, 2, 
/* out0093_had-eta15-phi12 */     0, 
/* out0094_had-eta15-phi13 */     1, 32, 2, 
/* out0095_had-eta15-phi14 */     1, 32, 2, 
/* out0096_had-eta16-phi12 */     0, 
/* out0097_had-eta16-phi13 */     0, 
/* out0098_had-eta12-phi15 */     2, 33, 2, 113, 2, 
/* out0099_had-eta12-phi16 */     2, 33, 2, 113, 2, 
/* out0100_had-eta12-phi17 */     2, 33, 2, 125, 2, 
/* out0101_had-eta13-phi15 */     3, 32, 2, 112, 2, 113, 2, 
/* out0102_had-eta13-phi16 */     1, 112, 2, 
/* out0103_had-eta13-phi17 */     1, 30, 2, 
/* out0104_had-eta14-phi15 */     2, 32, 2, 112, 2, 
/* out0105_had-eta14-phi16 */     2, 30, 2, 112, 2, 
/* out0106_had-eta9-phi17 */     1, 126, 4, 
/* out0107_had-eta9-phi18 */     0, 
/* out0108_had-eta10-phi16 */     2, 33, 2, 126, 2, 
/* out0109_had-eta10-phi17 */     2, 125, 2, 126, 2, 
/* out0110_had-eta10-phi18 */     1, 125, 2, 
/* out0111_had-eta11-phi17 */     2, 33, 2, 125, 4, 
/* out0112_had-eta11-phi18 */     2, 31, 2, 125, 4, 
/* out0113_had-eta7-phi18 */     0, 
/* out0114_had-eta7-phi19 */     0, 
/* out0115_had-eta8-phi18 */     0, 
/* out0116_had-eta8-phi19 */     0, 
/* out0117_had-eta5-phi19 */     0, 
/* out0118_had-eta5-phi20 */     0, 
/* out0119_had-eta6-phi19 */     0, 
/* out0120_had-eta6-phi20 */     1, 100, 2, 
/* out0121_had-eta4-phi19 */     0, 
/* out0122_had-eta4-phi20 */     1, 131, 6, 
/* out0123_had-eta2-phi20 */     2, 97, 2, 132, 1, 
/* out0124_had-eta3-phi20 */     2, 97, 4, 131, 2, 
/* out0125_had-eta1-phi20 */     1, 132, 2, 
/* out0126_had-eta1-phi21 */     1, 132, 2, 
/* out0127_had-eta0-phi21 */     1, 132, 2, 
/* out0128_had-eta0-phi22 */     3, 85, 2, 138, 2, 140, 2, 
/* out0129_had-eta12-phi1 */     0, 
/* out0130_had-eta12-phi2 */     0, 
/* out0131_had-eta13-phi1 */     0, 
/* out0132_had-eta13-phi2 */     0, 
/* out0133_had-eta13-phi3 */     0, 
/* out0134_had-eta14-phi1 */     0, 
/* out0135_had-eta14-phi2 */     0, 
/* out0136_had-eta14-phi3 */     0, 
/* out0137_had-eta13-phi4 */     0, 
/* out0138_had-eta13-phi5 */     0, 
/* out0139_had-eta13-phi6 */     0, 
/* out0140_had-eta13-phi7 */     0, 
/* out0141_had-eta14-phi4 */     0, 
/* out0142_had-eta14-phi5 */     0, 
/* out0143_had-eta14-phi6 */     0, 
/* out0144_had-eta14-phi7 */     0, 
/* out0145_had-eta12-phi9 */     0, 
/* out0146_had-eta12-phi10 */     0, 
/* out0147_had-eta13-phi8 */     0, 
/* out0148_had-eta13-phi9 */     0, 
/* out0149_had-eta13-phi10 */     0, 
/* out0150_had-eta14-phi8 */     0, 
/* out0151_had-eta14-phi9 */     0, 
/* out0152_had-eta14-phi10 */     0, 
/* out0153_had-eta11-phi12 */     1, 34, 2, 
/* out0154_had-eta11-phi13 */     1, 34, 2, 
/* out0155_had-eta12-phi11 */     0, 
/* out0156_had-eta12-phi12 */     0, 
/* out0157_had-eta12-phi13 */     1, 34, 2, 
/* out0158_had-eta12-phi14 */     1, 113, 2, 
/* out0159_had-eta13-phi12 */     0, 
/* out0160_had-eta13-phi13 */     1, 32, 2, 
/* out0161_had-eta9-phi14 */     1, 114, 4, 
/* out0162_had-eta9-phi15 */     1, 114, 2, 
/* out0163_had-eta9-phi16 */     1, 126, 4, 
/* out0164_had-eta10-phi14 */     2, 34, 2, 114, 4, 
/* out0165_had-eta10-phi15 */     2, 33, 2, 114, 2, 
/* out0166_had-eta11-phi14 */     2, 34, 2, 113, 2, 
/* out0167_had-eta11-phi15 */     2, 33, 2, 113, 4, 
/* out0168_had-eta7-phi16 */     2, 127, 6, 153, 2, 
/* out0169_had-eta7-phi17 */     1, 153, 2, 
/* out0170_had-eta8-phi15 */     1, 127, 2, 
/* out0171_had-eta8-phi16 */     3, 126, 2, 127, 4, 153, 2, 
/* out0172_had-eta8-phi17 */     2, 126, 2, 153, 2, 
/* out0173_had-eta5-phi17 */     3, 15, 6, 145, 3, 153, 1, 
/* out0174_had-eta5-phi18 */     1, 15, 6, 
/* out0175_had-eta6-phi17 */     3, 15, 2, 145, 1, 153, 3, 
/* out0176_had-eta6-phi18 */     1, 15, 2, 
/* out0177_had-eta4-phi18 */     0, 
/* out0178_had-eta2-phi19 */     1, 97, 4, 
/* out0179_had-eta3-phi18 */     1, 98, 10, 
/* out0180_had-eta3-phi19 */     2, 97, 6, 98, 2, 
/* out0181_had-eta1-phi19 */     0, 
/* out0182_had-eta0-phi20 */     1, 132, 2, 
/* out0183_had-eta9-phi1 */     2, 19, 2, 103, 2, 
/* out0184_had-eta9-phi2 */     2, 1, 2, 35, 2, 
/* out0185_had-eta10-phi0 */     0, 
/* out0186_had-eta10-phi1 */     0, 
/* out0187_had-eta10-phi2 */     0, 
/* out0188_had-eta11-phi0 */     0, 
/* out0189_had-eta11-phi1 */     0, 
/* out0190_had-eta11-phi2 */     0, 
/* out0191_had-eta10-phi3 */     0, 
/* out0192_had-eta10-phi4 */     1, 123, 2, 
/* out0193_had-eta10-phi5 */     2, 122, 2, 123, 2, 
/* out0194_had-eta11-phi3 */     0, 
/* out0195_had-eta11-phi4 */     0, 
/* out0196_had-eta11-phi5 */     1, 122, 4, 
/* out0197_had-eta12-phi4 */     0, 
/* out0198_had-eta12-phi5 */     1, 122, 2, 
/* out0199_had-eta10-phi6 */     1, 122, 2, 
/* out0200_had-eta10-phi7 */     0, 
/* out0201_had-eta10-phi8 */     0, 
/* out0202_had-eta11-phi6 */     1, 122, 4, 
/* out0203_had-eta11-phi7 */     0, 
/* out0204_had-eta11-phi8 */     0, 
/* out0205_had-eta12-phi7 */     0, 
/* out0206_had-eta12-phi8 */     0, 
/* out0207_had-eta9-phi9 */     0, 
/* out0208_had-eta9-phi10 */     1, 20, 2, 
/* out0209_had-eta10-phi9 */     0, 
/* out0210_had-eta10-phi10 */     0, 
/* out0211_had-eta10-phi11 */     0, 
/* out0212_had-eta11-phi9 */     0, 
/* out0213_had-eta11-phi10 */     0, 
/* out0214_had-eta11-phi11 */     0, 
/* out0215_had-eta8-phi12 */     1, 64, 2, 
/* out0216_had-eta8-phi13 */     1, 115, 2, 
/* out0217_had-eta9-phi11 */     0, 
/* out0218_had-eta9-phi12 */     0, 
/* out0219_had-eta9-phi13 */     2, 34, 2, 114, 2, 
/* out0220_had-eta10-phi12 */     1, 34, 2, 
/* out0221_had-eta7-phi13 */     2, 2, 2, 115, 4, 
/* out0222_had-eta7-phi14 */     1, 115, 6, 
/* out0223_had-eta7-phi15 */     1, 127, 4, 
/* out0224_had-eta8-phi14 */     2, 114, 2, 115, 4, 
/* out0225_had-eta5-phi15 */     0, 
/* out0226_had-eta5-phi16 */     2, 145, 3, 153, 1, 
/* out0227_had-eta6-phi15 */     0, 
/* out0228_had-eta6-phi16 */     2, 145, 1, 153, 3, 
/* out0229_had-eta4-phi16 */     3, 16, 4, 145, 4, 154, 1, 
/* out0230_had-eta4-phi17 */     3, 16, 6, 145, 4, 154, 1, 
/* out0231_had-eta3-phi17 */     3, 16, 4, 146, 1, 154, 1, 
/* out0232_had-eta1-phi18 */     0, 
/* out0233_had-eta2-phi18 */     1, 98, 4, 
/* out0234_had-eta0-phi19 */     0, 
/* out0235_had-eta7-phi0 */     6, 0, 2, 19, 2, 63, 4, 103, 2, 104, 4, 147, 2, 
/* out0236_had-eta7-phi1 */     6, 0, 4, 19, 2, 21, 2, 63, 2, 104, 2, 147, 2, 
/* out0237_had-eta7-phi2 */     5, 0, 2, 4, 2, 35, 4, 38, 2, 151, 2, 
/* out0238_had-eta8-phi0 */     5, 0, 2, 19, 4, 63, 4, 103, 4, 147, 2, 
/* out0239_had-eta8-phi1 */     6, 0, 4, 19, 4, 35, 2, 63, 2, 103, 2, 147, 2, 
/* out0240_had-eta8-phi2 */     5, 0, 2, 1, 2, 19, 2, 35, 4, 151, 2, 
/* out0241_had-eta7-phi3 */     6, 1, 2, 4, 2, 35, 2, 39, 4, 124, 4, 151, 2, 
/* out0242_had-eta8-phi3 */     5, 1, 4, 35, 2, 36, 2, 124, 2, 151, 2, 
/* out0243_had-eta8-phi4 */     4, 1, 2, 36, 4, 123, 2, 124, 2, 
/* out0244_had-eta9-phi3 */     1, 1, 2, 
/* out0245_had-eta9-phi4 */     3, 1, 2, 36, 2, 123, 4, 
/* out0246_had-eta8-phi5 */     2, 36, 4, 123, 2, 
/* out0247_had-eta8-phi6 */     3, 37, 4, 53, 2, 143, 2, 
/* out0248_had-eta9-phi5 */     2, 36, 2, 123, 4, 
/* out0249_had-eta9-phi6 */     1, 37, 2, 
/* out0250_had-eta7-phi8 */     3, 40, 4, 54, 4, 135, 2, 
/* out0251_had-eta8-phi7 */     3, 37, 4, 53, 2, 143, 2, 
/* out0252_had-eta8-phi8 */     2, 54, 2, 135, 2, 
/* out0253_had-eta8-phi9 */     3, 20, 2, 54, 2, 135, 2, 
/* out0254_had-eta9-phi7 */     1, 37, 4, 
/* out0255_had-eta9-phi8 */     0, 
/* out0256_had-eta7-phi9 */     2, 54, 4, 135, 2, 
/* out0257_had-eta7-phi10 */     4, 20, 2, 22, 2, 64, 2, 128, 8, 
/* out0258_had-eta7-phi11 */     4, 2, 2, 20, 2, 64, 4, 128, 8, 
/* out0259_had-eta8-phi10 */     2, 20, 4, 64, 2, 
/* out0260_had-eta8-phi11 */     2, 20, 4, 64, 4, 
/* out0261_had-eta6-phi11 */     3, 2, 2, 22, 4, 66, 4, 
/* out0262_had-eta6-phi12 */     2, 2, 4, 66, 2, 
/* out0263_had-eta6-phi13 */     2, 2, 2, 116, 6, 
/* out0264_had-eta7-phi12 */     2, 2, 4, 64, 2, 
/* out0265_had-eta5-phi13 */     3, 5, 2, 116, 4, 117, 4, 
/* out0266_had-eta5-phi14 */     2, 116, 2, 117, 2, 
/* out0267_had-eta6-phi14 */     1, 116, 4, 
/* out0268_had-eta4-phi14 */     1, 117, 2, 
/* out0269_had-eta4-phi15 */     0, 
/* out0270_had-eta2-phi16 */     4, 17, 8, 18, 2, 146, 1, 154, 2, 
/* out0271_had-eta3-phi15 */     0, 
/* out0272_had-eta3-phi16 */     4, 16, 2, 17, 6, 146, 1, 154, 1, 
/* out0273_had-eta1-phi17 */     2, 146, 1, 154, 2, 
/* out0274_had-eta2-phi17 */     3, 17, 2, 146, 1, 154, 2, 
/* out0275_had-eta5-phi0 */     7, 3, 4, 21, 2, 23, 2, 65, 6, 67, 2, 105, 8, 147, 2, 
/* out0276_had-eta5-phi1 */     9, 3, 4, 7, 2, 21, 2, 23, 2, 38, 2, 41, 2, 65, 2, 105, 2, 147, 2, 
/* out0277_had-eta6-phi0 */     5, 3, 4, 21, 4, 65, 4, 104, 6, 147, 2, 
/* out0278_had-eta6-phi1 */     6, 3, 4, 21, 6, 38, 4, 65, 2, 104, 2, 147, 2, 
/* out0279_had-eta5-phi2 */     6, 4, 2, 7, 4, 38, 2, 41, 2, 42, 2, 151, 2, 
/* out0280_had-eta6-phi2 */     3, 4, 6, 38, 6, 151, 2, 
/* out0281_had-eta6-phi3 */     3, 4, 4, 39, 4, 151, 2, 
/* out0282_had-eta6-phi4 */     3, 39, 4, 124, 2, 141, 2, 
/* out0283_had-eta6-phi5 */     1, 141, 2, 
/* out0284_had-eta7-phi4 */     3, 36, 2, 39, 4, 124, 6, 
/* out0285_had-eta7-phi5 */     0, 
/* out0286_had-eta6-phi6 */     3, 53, 2, 143, 2, 155, 3, 
/* out0287_had-eta6-phi7 */     5, 40, 4, 53, 2, 55, 4, 143, 2, 155, 3, 
/* out0288_had-eta7-phi6 */     2, 53, 4, 143, 2, 
/* out0289_had-eta7-phi7 */     4, 37, 2, 40, 4, 53, 4, 143, 2, 
/* out0290_had-eta5-phi8 */     5, 43, 6, 55, 4, 56, 2, 57, 2, 135, 2, 
/* out0291_had-eta5-phi9 */     3, 43, 2, 56, 8, 135, 2, 
/* out0292_had-eta6-phi8 */     4, 40, 4, 54, 2, 55, 2, 135, 2, 
/* out0293_had-eta6-phi9 */     3, 54, 2, 56, 2, 135, 2, 
/* out0294_had-eta5-phi10 */     4, 22, 2, 24, 2, 56, 2, 66, 2, 
/* out0295_had-eta5-phi11 */     5, 5, 2, 22, 2, 24, 2, 66, 6, 68, 2, 
/* out0296_had-eta6-phi10 */     2, 22, 6, 66, 2, 
/* out0297_had-eta4-phi12 */     3, 5, 4, 8, 4, 68, 2, 
/* out0298_had-eta4-phi13 */     2, 5, 2, 117, 8, 
/* out0299_had-eta5-phi12 */     1, 5, 6, 
/* out0300_had-eta3-phi13 */     1, 8, 2, 
/* out0301_had-eta3-phi14 */     0, 
/* out0302_had-eta2-phi14 */     0, 
/* out0303_had-eta2-phi15 */     1, 18, 2, 
/* out0304_had-eta1-phi15 */     1, 18, 4, 
/* out0305_had-eta1-phi16 */     3, 18, 8, 146, 1, 154, 2, 
/* out0306_had-eta0-phi16 */     2, 146, 2, 154, 2, 
/* out0307_had-eta3-phi0 */     7, 6, 2, 9, 4, 25, 6, 67, 2, 69, 8, 106, 8, 148, 1, 
/* out0308_had-eta3-phi1 */     6, 6, 2, 9, 2, 10, 4, 25, 4, 44, 8, 148, 1, 
/* out0309_had-eta4-phi0 */     6, 6, 6, 23, 6, 67, 8, 105, 4, 106, 6, 148, 1, 
/* out0310_had-eta4-phi1 */     6, 6, 6, 7, 2, 23, 6, 41, 8, 67, 2, 148, 1, 
/* out0311_had-eta4-phi2 */     7, 7, 6, 10, 2, 41, 4, 42, 2, 45, 2, 129, 8, 152, 1, 
/* out0312_had-eta4-phi3 */     5, 7, 2, 42, 4, 45, 2, 129, 8, 152, 1, 
/* out0313_had-eta4-phi4 */     1, 141, 2, 
/* out0314_had-eta5-phi3 */     2, 42, 6, 151, 2, 
/* out0315_had-eta5-phi4 */     2, 42, 2, 141, 4, 
/* out0316_had-eta4-phi5 */     1, 141, 2, 
/* out0317_had-eta4-phi6 */     2, 144, 1, 155, 1, 
/* out0318_had-eta5-phi5 */     1, 141, 4, 
/* out0319_had-eta5-phi6 */     2, 143, 2, 155, 4, 
/* out0320_had-eta4-phi7 */     3, 57, 4, 144, 1, 155, 1, 
/* out0321_had-eta4-phi8 */     4, 43, 4, 46, 2, 57, 8, 136, 1, 
/* out0322_had-eta5-phi7 */     4, 43, 2, 55, 6, 143, 2, 155, 4, 
/* out0323_had-eta4-phi9 */     5, 43, 2, 46, 2, 56, 2, 58, 6, 136, 1, 
/* out0324_had-eta4-phi10 */     3, 24, 6, 58, 4, 68, 2, 
/* out0325_had-eta3-phi10 */     3, 26, 4, 58, 2, 60, 2, 
/* out0326_had-eta3-phi11 */     4, 8, 2, 26, 8, 68, 2, 70, 8, 
/* out0327_had-eta4-phi11 */     2, 24, 6, 68, 8, 
/* out0328_had-eta3-phi12 */     2, 8, 8, 70, 2, 
/* out0329_had-eta2-phi13 */     1, 149, 5, 
/* out0330_had-eta1-phi14 */     0, 
/* out0331_had-eta0-phi15 */     0, 
/* out0332_had-eta2-phi0 */     8, 9, 6, 12, 2, 25, 4, 27, 6, 47, 2, 69, 6, 71, 4, 148, 1, 
/* out0333_had-eta2-phi1 */     7, 9, 4, 13, 6, 25, 2, 27, 2, 44, 4, 47, 8, 148, 1, 
/* out0334_had-eta2-phi2 */     6, 10, 2, 13, 4, 48, 10, 130, 1, 133, 4, 152, 1, 
/* out0335_had-eta3-phi2 */     5, 10, 8, 44, 4, 45, 6, 130, 1, 152, 1, 
/* out0336_had-eta3-phi3 */     3, 45, 6, 130, 1, 152, 1, 
/* out0337_had-eta3-phi4 */     1, 142, 1, 
/* out0338_had-eta3-phi5 */     1, 142, 1, 
/* out0339_had-eta3-phi6 */     3, 72, 8, 144, 1, 156, 1, 
/* out0340_had-eta3-phi7 */     3, 72, 2, 144, 1, 156, 1, 
/* out0341_had-eta3-phi8 */     4, 46, 6, 57, 2, 59, 6, 136, 1, 
/* out0342_had-eta2-phi9 */     5, 49, 10, 59, 2, 60, 6, 61, 4, 136, 1, 
/* out0343_had-eta3-phi9 */     5, 46, 6, 58, 4, 59, 4, 60, 2, 136, 1, 
/* out0344_had-eta2-phi10 */     4, 26, 2, 28, 2, 60, 6, 62, 2, 
/* out0345_had-eta2-phi11 */     5, 11, 2, 26, 2, 28, 6, 70, 6, 73, 6, 
/* out0346_had-eta1-phi12 */     4, 11, 4, 73, 2, 149, 3, 150, 1, 
/* out0347_had-eta2-phi12 */     2, 11, 10, 149, 5, 
/* out0348_had-eta1-phi13 */     2, 149, 3, 150, 1, 
/* out0349_had-eta0-phi13 */     1, 150, 5, 
/* out0350_had-eta0-phi14 */     0, 
/* out0351_had-eta1-phi0 */     5, 12, 10, 27, 6, 50, 2, 71, 10, 148, 2, 
/* out0352_had-eta1-phi1 */     8, 12, 4, 13, 4, 14, 6, 27, 2, 47, 6, 50, 8, 51, 2, 148, 2, 
/* out0353_had-eta1-phi2 */     7, 13, 2, 14, 2, 48, 2, 51, 12, 130, 2, 133, 4, 152, 2, 
/* out0354_had-eta2-phi3 */     4, 48, 4, 130, 1, 133, 4, 152, 1, 
/* out0355_had-eta2-phi4 */     1, 142, 1, 
/* out0356_had-eta2-phi5 */     3, 74, 4, 86, 8, 142, 1, 
/* out0357_had-eta2-phi6 */     6, 72, 4, 74, 6, 75, 2, 86, 8, 144, 1, 156, 1, 
/* out0358_had-eta2-phi7 */     4, 72, 2, 75, 6, 144, 1, 156, 1, 
/* out0359_had-eta2-phi8 */     4, 49, 4, 59, 4, 61, 2, 136, 1, 
/* out0360_had-eta1-phi9 */     6, 49, 2, 52, 12, 61, 6, 62, 4, 89, 2, 136, 2, 
/* out0361_had-eta1-phi10 */     3, 28, 2, 52, 2, 62, 10, 
/* out0362_had-eta1-phi11 */     2, 28, 6, 73, 8, 
/* out0363_had-eta0-phi1 */     3, 14, 6, 50, 4, 148, 2, 
/* out0364_had-eta0-phi2 */     5, 14, 2, 51, 2, 130, 2, 134, 7, 152, 2, 
/* out0365_had-eta1-phi3 */     3, 130, 2, 133, 4, 152, 2, 
/* out0366_had-eta1-phi4 */     3, 76, 2, 87, 2, 142, 1, 
/* out0367_had-eta1-phi5 */     4, 74, 2, 76, 10, 87, 14, 142, 1, 
/* out0368_had-eta1-phi6 */     5, 74, 4, 75, 2, 88, 14, 144, 2, 156, 2, 
/* out0369_had-eta1-phi7 */     4, 75, 6, 88, 2, 144, 2, 156, 2, 
/* out0370_had-eta1-phi8 */     3, 61, 4, 89, 8, 136, 2, 
/* out0371_had-eta0-phi9 */     4, 52, 2, 89, 2, 93, 10, 136, 2, 
/* out0372_had-eta0-phi10 */     0, 
/* out0373_had-eta16-phi20 */     0, 
/* out0374_had-eta16-phi21 */     1, 77, 2, 
/* out0375_had-eta17-phi19 */     0, 
/* out0376_had-eta17-phi20 */     0, 
/* out0377_had-eta17-phi21 */     0, 
/* out0378_had-eta17-phi22 */     1, 77, 2, 
/* out0379_had-eta12-phi21 */     1, 95, 2, 
/* out0380_had-eta13-phi21 */     0, 
/* out0381_had-eta14-phi20 */     1, 94, 2, 
/* out0382_had-eta11-phi21 */     1, 95, 2, 
/* out0383_had-eta16-phi14 */     1, 29, 2, 
/* out0384_had-eta16-phi15 */     1, 29, 2, 
/* out0385_had-eta17-phi13 */     1, 29, 2, 
/* out0386_had-eta17-phi14 */     1, 29, 2, 
/* out0387_had-eta17-phi15 */     1, 29, 2, 
/* out0388_had-eta17-phi16 */     1, 29, 2, 
/* out0389_had-eta17-phi17 */     1, 29, 2, 
/* out0390_had-eta14-phi17 */     2, 30, 2, 112, 2, 
/* out0391_had-eta14-phi18 */     2, 30, 2, 94, 2, 
/* out0392_had-eta14-phi0 */     0, 
/* out0393_had-eta15-phi0 */     0, 
/* out0394_had-eta15-phi1 */     0, 
/* out0395_had-eta15-phi2 */     0, 
/* out0396_had-eta16-phi0 */     0, 
/* out0397_had-eta15-phi4 */     0, 
/* out0398_had-eta15-phi5 */     0, 
/* out0399_had-eta15-phi6 */     0, 
/* out0400_had-eta16-phi5 */     0, 
/* out0401_had-eta16-phi6 */     0, 
/* out0402_had-eta14-phi11 */     0, 
/* out0403_had-eta15-phi9 */     0, 
/* out0404_had-eta15-phi10 */     0, 
/* out0405_had-eta15-phi11 */     0, 
/* out0406_had-eta16-phi11 */     0, 
/* out0407_had-eta13-phi14 */     1, 32, 2, 
/* out0408_had-eta11-phi16 */     2, 33, 2, 113, 2, 
/* out0409_had-eta12-phi-1 */     0, 
/* out0410_had-eta12-phi0 */     0, 
/* out0411_had-eta13-phi0 */     0, 
/* out0412_had-eta12-phi3 */     0, 
/* out0413_had-eta12-phi6 */     1, 122, 2, 
/* out0414_had-eta13-phi11 */     0, 
/* out0415_had-eta10-phi13 */     1, 34, 2, 
/* out0416_had-eta9-phi-1 */     0, 
/* out0417_had-eta9-phi0 */     1, 103, 4, 
/* out0418_had-eta0-phi18 */     0, 
/* out0419_had-eta7-phi-1 */     1, 63, 2, 
/* out0420_had-eta5-phi-1 */     2, 65, 2, 105, 2, 
/* out0421_had-eta0-phi17 */     2, 146, 2, 154, 2, 
/* out0422_had-eta3-phi-1 */     2, 69, 2, 106, 2, 
/* out0423_had-eta2-phi-1 */     0, 
/* out0424_had-eta0-phi0 */     2, 50, 2, 148, 2, 
/* out0425_had-eta1-phi-1 */     1, 71, 2, 
/* out0426_had-eta0-phi11 */     0, 
/* out0427_had-eta0-phi3 */     3, 130, 2, 134, 7, 152, 2, 
/* out0428_had-eta0-phi8 */     4, 89, 4, 92, 10, 93, 6, 136, 2, 
/* out0429_had-eta16-phi23 */     1, 77, 2, 
/* out0430_had-eta4-phi24 */     0, 
/* out0431_had-eta0-phi23 */     3, 85, 14, 138, 2, 140, 2, 
/* out0432_had-eta1-phi24 */     0, 
/* out0433_had-eta17-phi5 */     0, 
/* out0434_had-eta17-phi7 */     0, 
/* out0435_had-eta0-phi12 */     1, 150, 5, 
/* out0436_had-eta0-phi4 */     2, 90, 8, 142, 2, 
/* out0437_had-eta0-phi5 */     3, 76, 4, 90, 8, 142, 2, 
/* out0438_had-eta0-phi6 */     3, 91, 8, 144, 2, 156, 2, 
/* out0439_had-eta0-phi7 */     4, 91, 8, 92, 6, 144, 2, 156, 2, 
/* out0440_had-eta17-phi18 */     0, 
/* out0441_had-eta16-phi-1 */     0, 
/* out0442_had-eta17-phi11 */     0, 
/* out0443_had-eta4-phi-1 */     1, 67, 2, 
/* out0444_had-eta16-phi24 */     0, 
/* out0445_had-eta17-phi23 */     1, 77, 2, 
/* out0446_had-eta10-phi24 */     1, 79, 2, 
/* out0447_had-eta17-phi12 */     0, 
/* out0448_had-eta15-phi7 */     0, 
/* out0449_had-eta17-phi0 */     0, 
/* out0450_had-eta15-phi15 */     1, 112, 2, 
/* out0451_had-eta10-phi-1 */     0, 
/* out0452_had-eta8-phi-1 */     2, 63, 2, 103, 2, 
/* out0453_had-eta13-phi24 */     2, 78, 2, 107, 2, 
/* out0454_had-eta8-phi24 */     1, 109, 2, 
/* out0455_had-eta0-phi24 */     0, 
/* out0456_had-eta15-phi8 */     0, 
/* out0457_had-eta13-phi-1 */     0, 
/* out0458_had-eta15-phi3 */     0, 
/* out0459_had-eta6-phi-1 */     1, 104, 2, 
/* out0460_had-eta15-phi20 */     1, 94, 2, 
/* out0461_had-eta17-phi24 */     0, 
/* out0462_had-eta17-phi-1 */     0, 
/* out0463_had-eta11-phi-1 */     0, 
/* out0464_had-eta14-phi24 */     2, 107, 2, 118, 2, 
/* out0465_had-eta14-phi-1 */     0, 
/* out0466_had-eta15-phi-1 */     0, 
/* out0467_had-eta-2-phi0 */     0, 
/* out0468_had-eta-1-phi0 */     1, 148, 1, 
/* out0469_had-eta-2-phi1 */     0, 
/* out0470_had-eta-1-phi1 */     1, 148, 1, 
/* out0471_had-eta-2-phi2 */     0, 
/* out0472_had-eta-1-phi2 */     3, 130, 2, 134, 1, 152, 1, 
/* out0473_had-eta-2-phi3 */     0, 
/* out0474_had-eta-1-phi3 */     3, 130, 2, 134, 1, 152, 1, 
/* out0475_had-eta-2-phi4 */     1, 142, 1, 
/* out0476_had-eta-1-phi4 */     1, 142, 2, 
/* out0477_had-eta-2-phi5 */     1, 142, 1, 
/* out0478_had-eta-1-phi5 */     1, 142, 2, 
/* out0479_had-eta-2-phi6 */     0, 
/* out0480_had-eta-1-phi6 */     2, 144, 1, 156, 2, 
/* out0481_had-eta-2-phi7 */     0, 
/* out0482_had-eta-1-phi7 */     2, 144, 1, 156, 2, 
/* out0483_had-eta-2-phi8 */     0, 
/* out0484_had-eta-1-phi8 */     1, 136, 1, 
/* out0485_had-eta-2-phi9 */     0, 
/* out0486_had-eta-1-phi9 */     1, 136, 1, 
/* out0487_had-eta-2-phi10 */     0, 
/* out0488_had-eta-1-phi10 */     0, 
/* out0489_had-eta-2-phi11 */     0, 
/* out0490_had-eta-1-phi11 */     0, 
/* out0491_had-eta-2-phi12 */     0, 
/* out0492_had-eta-1-phi12 */     1, 150, 2, 
/* out0493_had-eta-2-phi13 */     0, 
/* out0494_had-eta-1-phi13 */     1, 150, 2, 
/* out0495_had-eta-2-phi14 */     0, 
/* out0496_had-eta-1-phi14 */     0, 
/* out0497_had-eta-2-phi15 */     0, 
/* out0498_had-eta-1-phi15 */     0, 
/* out0499_had-eta-2-phi16 */     1, 146, 1, 
/* out0500_had-eta-1-phi16 */     1, 146, 2, 
/* out0501_had-eta-2-phi17 */     1, 146, 1, 
/* out0502_had-eta-1-phi17 */     1, 146, 2, 
/* out0503_had-eta-2-phi18 */     0, 
/* out0504_had-eta-1-phi18 */     0, 
/* out0505_had-eta-2-phi19 */     0, 
/* out0506_had-eta-1-phi19 */     0, 
/* out0507_had-eta-2-phi20 */     0, 
/* out0508_had-eta-1-phi20 */     1, 132, 3, 
/* out0509_had-eta-2-phi21 */     0, 
/* out0510_had-eta-1-phi21 */     1, 132, 3, 
/* out0511_had-eta-2-phi22 */     0, 
/* out0512_had-eta-1-phi22 */     1, 140, 2, 
/* out0513_had-eta-2-phi23 */     0, 
/* out0514_had-eta-1-phi23 */     11402
};