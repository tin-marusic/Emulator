parameter integer matrixE [0:1437] = {
/* num inputs = 106 (in0-in105) */
/* num outputs = 428(out0-out427) */
//* max inputs per outputs = 5 */
//* total number of input in adders 505 */

/* out0000_em-eta16-phi16 */     0, 
/* out0001_em-eta16-phi17 */     0, 
/* out0002_em-eta16-phi18 */     0, 
/* out0003_em-eta16-phi19 */     0, 
/* out0004_em-eta17-phi15 */     0, 
/* out0005_em-eta17-phi16 */     0, 
/* out0006_em-eta17-phi17 */     1, 81, 1, 
/* out0007_em-eta17-phi18 */     1, 81, 1, 
/* out0008_em-eta12-phi19 */     0, 
/* out0009_em-eta12-phi20 */     1, 83, 1, 
/* out0010_em-eta12-phi21 */     1, 83, 1, 
/* out0011_em-eta13-phi18 */     0, 
/* out0012_em-eta13-phi19 */     1, 82, 1, 
/* out0013_em-eta13-phi20 */     1, 82, 1, 
/* out0014_em-eta13-phi21 */     0, 
/* out0015_em-eta14-phi20 */     1, 82, 1, 
/* out0016_em-eta9-phi20 */     1, 50, 1, 
/* out0017_em-eta9-phi21 */     0, 
/* out0018_em-eta9-phi22 */     0, 
/* out0019_em-eta10-phi20 */     1, 83, 1, 
/* out0020_em-eta10-phi21 */     1, 83, 1, 
/* out0021_em-eta10-phi22 */     1, 83, 1, 
/* out0022_em-eta11-phi20 */     1, 83, 1, 
/* out0023_em-eta11-phi21 */     1, 83, 1, 
/* out0024_em-eta6-phi21 */     3, 52, 1, 73, 2, 84, 2, 
/* out0025_em-eta6-phi22 */     2, 73, 2, 84, 2, 
/* out0026_em-eta7-phi20 */     1, 52, 2, 
/* out0027_em-eta7-phi21 */     1, 84, 1, 
/* out0028_em-eta7-phi22 */     2, 73, 1, 84, 1, 
/* out0029_em-eta8-phi21 */     0, 
/* out0030_em-eta8-phi22 */     0, 
/* out0031_em-eta4-phi21 */     4, 53, 2, 54, 1, 74, 1, 85, 1, 
/* out0032_em-eta4-phi22 */     2, 74, 3, 85, 3, 
/* out0033_em-eta5-phi21 */     3, 53, 1, 73, 1, 85, 1, 
/* out0034_em-eta5-phi22 */     4, 73, 1, 74, 2, 84, 1, 85, 2, 
/* out0035_em-eta5-phi23 */     0, 
/* out0036_em-eta2-phi22 */     5, 55, 1, 75, 3, 76, 1, 86, 2, 87, 2, 
/* out0037_em-eta3-phi21 */     1, 54, 4, 
/* out0038_em-eta3-phi22 */     3, 74, 1, 75, 3, 86, 4, 
/* out0039_em-eta3-phi23 */     2, 75, 1, 86, 2, 
/* out0040_em-eta1-phi22 */     4, 55, 1, 56, 1, 76, 4, 87, 3, 
/* out0041_em-eta1-phi23 */     2, 76, 2, 87, 2, 
/* out0042_em-eta2-phi23 */     3, 75, 1, 76, 1, 87, 1, 
/* out0043_em-eta0-phi22 */     1, 56, 2, 
/* out0044_em-eta0-phi23 */     0, 
/* out0045_em-eta15-phi-2 */     0, 
/* out0046_em-eta15-phi-1 */     0, 
/* out0047_em-eta15-phi0 */     0, 
/* out0048_em-eta15-phi1 */     0, 
/* out0049_em-eta16-phi-3 */     0, 
/* out0050_em-eta16-phi-1 */     0, 
/* out0051_em-eta16-phi0 */     0, 
/* out0052_em-eta16-phi2 */     0, 
/* out0053_em-eta16-phi4 */     0, 
/* out0054_em-eta16-phi5 */     1, 13, 1, 
/* out0055_em-eta16-phi6 */     1, 13, 1, 
/* out0056_em-eta16-phi7 */     0, 
/* out0057_em-eta17-phi5 */     2, 13, 1, 65, 1, 
/* out0058_em-eta17-phi6 */     2, 13, 1, 65, 1, 
/* out0059_em-eta17-phi7 */     2, 13, 1, 65, 1, 
/* out0060_em-eta17-phi8 */     0, 
/* out0061_em-eta15-phi10 */     0, 
/* out0062_em-eta15-phi11 */     0, 
/* out0063_em-eta15-phi12 */     0, 
/* out0064_em-eta15-phi13 */     0, 
/* out0065_em-eta16-phi10 */     1, 66, 1, 
/* out0066_em-eta16-phi12 */     1, 66, 1, 
/* out0067_em-eta16-phi13 */     1, 66, 1, 
/* out0068_em-eta17-phi12 */     1, 66, 1, 
/* out0069_em-eta12-phi14 */     0, 
/* out0070_em-eta12-phi15 */     1, 8, 1, 
/* out0071_em-eta12-phi16 */     1, 8, 1, 
/* out0072_em-eta13-phi14 */     1, 8, 1, 
/* out0073_em-eta13-phi15 */     1, 8, 1, 
/* out0074_em-eta13-phi16 */     1, 8, 1, 
/* out0075_em-eta13-phi17 */     1, 8, 1, 
/* out0076_em-eta14-phi16 */     0, 
/* out0077_em-eta9-phi17 */     1, 51, 1, 
/* out0078_em-eta9-phi18 */     1, 50, 1, 
/* out0079_em-eta10-phi16 */     0, 
/* out0080_em-eta10-phi17 */     1, 49, 1, 
/* out0081_em-eta10-phi18 */     1, 49, 1, 
/* out0082_em-eta10-phi19 */     0, 
/* out0083_em-eta11-phi17 */     1, 49, 1, 
/* out0084_em-eta11-phi18 */     1, 49, 1, 
/* out0085_em-eta7-phi18 */     1, 88, 2, 
/* out0086_em-eta7-phi19 */     2, 50, 1, 52, 1, 
/* out0087_em-eta8-phi18 */     2, 50, 1, 88, 1, 
/* out0088_em-eta8-phi19 */     1, 50, 2, 
/* out0089_em-eta8-phi20 */     1, 50, 1, 
/* out0090_em-eta9-phi19 */     1, 50, 1, 
/* out0091_em-eta5-phi19 */     1, 89, 2, 
/* out0092_em-eta5-phi20 */     1, 53, 2, 
/* out0093_em-eta6-phi19 */     2, 52, 2, 89, 1, 
/* out0094_em-eta6-phi20 */     1, 52, 2, 
/* out0095_em-eta3-phi20 */     4, 15, 1, 54, 2, 90, 1, 91, 1, 
/* out0096_em-eta4-phi20 */     2, 53, 3, 90, 1, 
/* out0097_em-eta2-phi20 */     4, 15, 1, 16, 2, 91, 4, 92, 1, 
/* out0098_em-eta2-phi21 */     2, 54, 1, 55, 3, 
/* out0099_em-eta0-phi21 */     2, 17, 1, 56, 3, 
/* out0100_em-eta1-phi21 */     3, 55, 3, 56, 2, 92, 1, 
/* out0101_em-eta11-phi-1 */     0, 
/* out0102_em-eta11-phi0 */     0, 
/* out0103_em-eta11-phi1 */     2, 18, 1, 43, 1, 
/* out0104_em-eta12-phi-2 */     0, 
/* out0105_em-eta12-phi-1 */     0, 
/* out0106_em-eta12-phi0 */     0, 
/* out0107_em-eta12-phi1 */     0, 
/* out0108_em-eta13-phi0 */     0, 
/* out0109_em-eta12-phi2 */     1, 43, 1, 
/* out0110_em-eta12-phi3 */     1, 14, 1, 
/* out0111_em-eta12-phi4 */     1, 14, 1, 
/* out0112_em-eta13-phi2 */     2, 14, 1, 42, 1, 
/* out0113_em-eta13-phi3 */     2, 14, 1, 42, 1, 
/* out0114_em-eta13-phi4 */     2, 14, 1, 42, 1, 
/* out0115_em-eta13-phi5 */     2, 14, 1, 42, 1, 
/* out0116_em-eta14-phi3 */     1, 42, 1, 
/* out0117_em-eta12-phi7 */     0, 
/* out0118_em-eta12-phi8 */     0, 
/* out0119_em-eta12-phi9 */     0, 
/* out0120_em-eta13-phi6 */     0, 
/* out0121_em-eta13-phi7 */     1, 67, 1, 
/* out0122_em-eta13-phi8 */     1, 67, 1, 
/* out0123_em-eta13-phi9 */     1, 67, 1, 
/* out0124_em-eta14-phi7 */     1, 67, 1, 
/* out0125_em-eta11-phi11 */     0, 
/* out0126_em-eta11-phi12 */     0, 
/* out0127_em-eta12-phi10 */     0, 
/* out0128_em-eta12-phi11 */     1, 68, 1, 
/* out0129_em-eta12-phi12 */     1, 68, 1, 
/* out0130_em-eta12-phi13 */     1, 68, 1, 
/* out0131_em-eta13-phi11 */     1, 68, 1, 
/* out0132_em-eta13-phi12 */     1, 68, 1, 
/* out0133_em-eta9-phi13 */     1, 9, 1, 
/* out0134_em-eta9-phi14 */     1, 9, 1, 
/* out0135_em-eta9-phi15 */     2, 9, 1, 51, 1, 
/* out0136_em-eta10-phi13 */     1, 9, 1, 
/* out0137_em-eta10-phi14 */     1, 9, 1, 
/* out0138_em-eta10-phi15 */     1, 9, 1, 
/* out0139_em-eta11-phi14 */     1, 9, 1, 
/* out0140_em-eta11-phi15 */     1, 9, 1, 
/* out0141_em-eta7-phi15 */     3, 10, 1, 57, 2, 101, 2, 
/* out0142_em-eta7-phi16 */     3, 51, 1, 57, 1, 101, 2, 
/* out0143_em-eta7-phi17 */     1, 88, 2, 
/* out0144_em-eta8-phi15 */     2, 51, 1, 101, 1, 
/* out0145_em-eta8-phi16 */     1, 51, 2, 
/* out0146_em-eta8-phi17 */     2, 51, 1, 88, 1, 
/* out0147_em-eta9-phi16 */     1, 51, 1, 
/* out0148_em-eta5-phi17 */     2, 0, 1, 93, 3, 
/* out0149_em-eta5-phi18 */     1, 89, 3, 
/* out0150_em-eta6-phi17 */     2, 88, 1, 93, 1, 
/* out0151_em-eta6-phi18 */     2, 88, 1, 89, 1, 
/* out0152_em-eta3-phi18 */     1, 23, 3, 
/* out0153_em-eta3-phi19 */     3, 15, 4, 90, 3, 91, 1, 
/* out0154_em-eta4-phi18 */     1, 89, 1, 
/* out0155_em-eta4-phi19 */     1, 90, 3, 
/* out0156_em-eta2-phi19 */     4, 15, 2, 16, 1, 24, 1, 91, 2, 
/* out0157_em-eta1-phi19 */     3, 16, 2, 24, 1, 25, 3, 
/* out0158_em-eta1-phi20 */     3, 16, 3, 17, 2, 92, 6, 
/* out0159_em-eta0-phi20 */     1, 17, 5, 
/* out0160_em-eta8-phi-1 */     0, 
/* out0161_em-eta8-phi0 */     0, 
/* out0162_em-eta9-phi-1 */     0, 
/* out0163_em-eta9-phi0 */     0, 
/* out0164_em-eta9-phi1 */     0, 
/* out0165_em-eta10-phi-1 */     0, 
/* out0166_em-eta10-phi0 */     0, 
/* out0167_em-eta9-phi2 */     3, 18, 1, 43, 1, 44, 1, 
/* out0168_em-eta9-phi3 */     2, 18, 1, 40, 1, 
/* out0169_em-eta10-phi1 */     2, 18, 1, 43, 1, 
/* out0170_em-eta10-phi2 */     2, 18, 1, 43, 1, 
/* out0171_em-eta10-phi3 */     2, 18, 1, 43, 1, 
/* out0172_em-eta11-phi2 */     2, 18, 1, 43, 1, 
/* out0173_em-eta11-phi3 */     2, 18, 1, 43, 1, 
/* out0174_em-eta9-phi5 */     1, 40, 1, 
/* out0175_em-eta9-phi6 */     1, 41, 1, 
/* out0176_em-eta10-phi4 */     0, 
/* out0177_em-eta10-phi5 */     1, 39, 1, 
/* out0178_em-eta10-phi6 */     1, 39, 1, 
/* out0179_em-eta10-phi7 */     0, 
/* out0180_em-eta11-phi5 */     1, 39, 1, 
/* out0181_em-eta11-phi6 */     1, 39, 1, 
/* out0182_em-eta9-phi8 */     1, 41, 1, 
/* out0183_em-eta9-phi9 */     0, 
/* out0184_em-eta9-phi10 */     0, 
/* out0185_em-eta10-phi8 */     0, 
/* out0186_em-eta10-phi9 */     0, 
/* out0187_em-eta10-phi10 */     0, 
/* out0188_em-eta11-phi8 */     0, 
/* out0189_em-eta11-phi9 */     0, 
/* out0190_em-eta8-phi11 */     0, 
/* out0191_em-eta8-phi12 */     0, 
/* out0192_em-eta9-phi11 */     0, 
/* out0193_em-eta9-phi12 */     0, 
/* out0194_em-eta10-phi11 */     0, 
/* out0195_em-eta10-phi12 */     0, 
/* out0196_em-eta6-phi13 */     1, 11, 1, 
/* out0197_em-eta6-phi14 */     2, 10, 1, 11, 1, 
/* out0198_em-eta7-phi13 */     1, 10, 2, 
/* out0199_em-eta7-phi14 */     1, 10, 2, 
/* out0200_em-eta8-phi13 */     1, 10, 1, 
/* out0201_em-eta8-phi14 */     1, 10, 1, 
/* out0202_em-eta5-phi15 */     3, 57, 1, 58, 2, 102, 3, 
/* out0203_em-eta5-phi16 */     1, 93, 2, 
/* out0204_em-eta6-phi15 */     3, 57, 2, 101, 2, 102, 1, 
/* out0205_em-eta6-phi16 */     3, 57, 2, 93, 1, 101, 1, 
/* out0206_em-eta3-phi16 */     4, 0, 1, 1, 3, 94, 2, 95, 1, 
/* out0207_em-eta3-phi17 */     2, 0, 1, 23, 3, 
/* out0208_em-eta4-phi16 */     3, 0, 2, 93, 1, 94, 3, 
/* out0209_em-eta4-phi17 */     2, 0, 3, 94, 1, 
/* out0210_em-eta2-phi17 */     2, 23, 1, 27, 4, 
/* out0211_em-eta2-phi18 */     2, 23, 1, 24, 4, 
/* out0212_em-eta1-phi18 */     3, 24, 2, 25, 1, 28, 2, 
/* out0213_em-eta0-phi18 */     2, 25, 1, 28, 2, 
/* out0214_em-eta0-phi19 */     1, 25, 3, 
/* out0215_em-eta5-phi-1 */     1, 29, 2, 
/* out0216_em-eta5-phi0 */     1, 29, 2, 
/* out0217_em-eta6-phi-1 */     1, 26, 2, 
/* out0218_em-eta6-phi0 */     1, 26, 2, 
/* out0219_em-eta7-phi-1 */     1, 26, 2, 
/* out0220_em-eta7-phi0 */     1, 26, 2, 
/* out0221_em-eta6-phi1 */     0, 
/* out0222_em-eta6-phi2 */     0, 
/* out0223_em-eta7-phi1 */     2, 19, 2, 44, 1, 
/* out0224_em-eta7-phi2 */     2, 19, 2, 44, 2, 
/* out0225_em-eta7-phi3 */     1, 19, 1, 
/* out0226_em-eta8-phi1 */     2, 19, 1, 44, 1, 
/* out0227_em-eta8-phi2 */     2, 19, 2, 44, 2, 
/* out0228_em-eta7-phi4 */     1, 40, 1, 
/* out0229_em-eta7-phi5 */     0, 
/* out0230_em-eta8-phi3 */     2, 40, 1, 44, 1, 
/* out0231_em-eta8-phi4 */     1, 40, 2, 
/* out0232_em-eta8-phi5 */     1, 40, 1, 
/* out0233_em-eta9-phi4 */     1, 40, 1, 
/* out0234_em-eta7-phi6 */     0, 
/* out0235_em-eta7-phi7 */     2, 30, 1, 41, 1, 
/* out0236_em-eta7-phi8 */     1, 30, 1, 
/* out0237_em-eta8-phi6 */     1, 41, 1, 
/* out0238_em-eta8-phi7 */     1, 41, 2, 
/* out0239_em-eta8-phi8 */     1, 41, 1, 
/* out0240_em-eta9-phi7 */     1, 41, 1, 
/* out0241_em-eta6-phi9 */     1, 69, 2, 
/* out0242_em-eta6-phi10 */     1, 69, 2, 
/* out0243_em-eta7-phi9 */     0, 
/* out0244_em-eta7-phi10 */     1, 69, 1, 
/* out0245_em-eta8-phi9 */     0, 
/* out0246_em-eta8-phi10 */     0, 
/* out0247_em-eta5-phi11 */     0, 
/* out0248_em-eta5-phi12 */     1, 11, 1, 
/* out0249_em-eta6-phi11 */     0, 
/* out0250_em-eta6-phi12 */     0, 
/* out0251_em-eta7-phi11 */     0, 
/* out0252_em-eta7-phi12 */     0, 
/* out0253_em-eta4-phi13 */     2, 11, 1, 12, 2, 
/* out0254_em-eta4-phi14 */     5, 12, 1, 58, 2, 59, 1, 102, 1, 103, 2, 
/* out0255_em-eta5-phi13 */     1, 11, 2, 
/* out0256_em-eta5-phi14 */     3, 11, 2, 58, 1, 102, 2, 
/* out0257_em-eta3-phi14 */     4, 12, 1, 59, 4, 103, 3, 104, 1, 
/* out0258_em-eta3-phi15 */     5, 1, 1, 59, 2, 94, 1, 95, 1, 103, 2, 
/* out0259_em-eta4-phi15 */     4, 58, 3, 94, 1, 102, 1, 103, 1, 
/* out0260_em-eta2-phi15 */     4, 1, 1, 2, 1, 95, 4, 96, 1, 
/* out0261_em-eta2-phi16 */     3, 1, 3, 27, 1, 95, 2, 
/* out0262_em-eta1-phi16 */     3, 2, 3, 27, 1, 31, 3, 
/* out0263_em-eta1-phi17 */     3, 27, 2, 28, 2, 31, 1, 
/* out0264_em-eta0-phi17 */     2, 28, 2, 31, 1, 
/* out0265_em-eta3-phi0 */     1, 32, 3, 
/* out0266_em-eta4-phi-1 */     1, 29, 2, 
/* out0267_em-eta4-phi0 */     1, 29, 2, 
/* out0268_em-eta4-phi1 */     0, 
/* out0269_em-eta4-phi2 */     1, 5, 2, 
/* out0270_em-eta5-phi1 */     0, 
/* out0271_em-eta5-phi2 */     0, 
/* out0272_em-eta5-phi3 */     1, 4, 2, 
/* out0273_em-eta5-phi4 */     3, 4, 2, 45, 2, 77, 2, 
/* out0274_em-eta6-phi3 */     1, 4, 2, 
/* out0275_em-eta6-phi4 */     1, 4, 2, 
/* out0276_em-eta5-phi5 */     2, 45, 2, 77, 3, 
/* out0277_em-eta5-phi6 */     0, 
/* out0278_em-eta6-phi5 */     1, 77, 1, 
/* out0279_em-eta6-phi6 */     0, 
/* out0280_em-eta5-phi7 */     1, 30, 1, 
/* out0281_em-eta5-phi8 */     2, 30, 1, 33, 1, 
/* out0282_em-eta6-phi7 */     1, 30, 2, 
/* out0283_em-eta6-phi8 */     1, 30, 2, 
/* out0284_em-eta4-phi9 */     2, 33, 2, 70, 1, 
/* out0285_em-eta4-phi10 */     1, 70, 4, 
/* out0286_em-eta5-phi9 */     2, 33, 1, 69, 1, 
/* out0287_em-eta5-phi10 */     2, 69, 2, 70, 1, 
/* out0288_em-eta3-phi12 */     1, 12, 1, 
/* out0289_em-eta4-phi11 */     1, 70, 1, 
/* out0290_em-eta4-phi12 */     0, 
/* out0291_em-eta2-phi13 */     2, 60, 1, 104, 1, 
/* out0292_em-eta3-phi13 */     1, 12, 3, 
/* out0293_em-eta2-phi14 */     3, 59, 1, 60, 3, 104, 5, 
/* out0294_em-eta1-phi15 */     2, 2, 4, 96, 6, 
/* out0295_em-eta0-phi16 */     1, 31, 3, 
/* out0296_em-eta2-phi-1 */     2, 32, 1, 34, 2, 
/* out0297_em-eta2-phi0 */     2, 32, 1, 34, 2, 
/* out0298_em-eta3-phi-1 */     1, 32, 3, 
/* out0299_em-eta2-phi1 */     0, 
/* out0300_em-eta3-phi1 */     0, 
/* out0301_em-eta3-phi2 */     2, 5, 1, 6, 1, 
/* out0302_em-eta3-phi3 */     5, 5, 2, 6, 1, 46, 2, 78, 1, 79, 1, 
/* out0303_em-eta4-phi3 */     2, 5, 3, 78, 1, 
/* out0304_em-eta3-phi4 */     2, 46, 4, 78, 3, 
/* out0305_em-eta3-phi5 */     3, 61, 2, 78, 1, 97, 1, 
/* out0306_em-eta4-phi4 */     4, 45, 2, 46, 1, 77, 1, 78, 2, 
/* out0307_em-eta4-phi5 */     4, 45, 2, 61, 1, 77, 1, 97, 2, 
/* out0308_em-eta3-phi6 */     4, 61, 3, 63, 1, 97, 2, 98, 3, 
/* out0309_em-eta3-phi7 */     1, 98, 1, 
/* out0310_em-eta4-phi6 */     2, 61, 2, 97, 3, 
/* out0311_em-eta4-phi7 */     0, 
/* out0312_em-eta3-phi8 */     2, 33, 1, 35, 1, 
/* out0313_em-eta3-phi9 */     1, 35, 3, 
/* out0314_em-eta4-phi8 */     1, 33, 3, 
/* out0315_em-eta2-phi10 */     2, 71, 3, 72, 1, 
/* out0316_em-eta3-phi10 */     2, 70, 1, 71, 3, 
/* out0317_em-eta3-phi11 */     1, 71, 1, 
/* out0318_em-eta2-phi11 */     2, 71, 1, 72, 1, 
/* out0319_em-eta2-phi12 */     0, 
/* out0320_em-eta1-phi12 */     0, 
/* out0321_em-eta1-phi13 */     3, 60, 1, 62, 1, 105, 2, 
/* out0322_em-eta0-phi14 */     3, 3, 1, 62, 3, 105, 1, 
/* out0323_em-eta1-phi14 */     5, 60, 3, 62, 2, 96, 1, 104, 1, 105, 4, 
/* out0324_em-eta0-phi15 */     1, 3, 7, 
/* out0325_em-eta1-phi-1 */     2, 34, 2, 36, 1, 
/* out0326_em-eta1-phi0 */     2, 34, 2, 36, 1, 
/* out0327_em-eta1-phi1 */     1, 7, 1, 
/* out0328_em-eta2-phi2 */     1, 6, 4, 
/* out0329_em-eta2-phi3 */     3, 6, 2, 47, 3, 79, 4, 
/* out0330_em-eta2-phi4 */     3, 46, 1, 47, 2, 79, 3, 
/* out0331_em-eta2-phi5 */     0, 
/* out0332_em-eta2-phi6 */     3, 20, 3, 63, 5, 98, 3, 
/* out0333_em-eta2-phi7 */     4, 20, 1, 63, 2, 98, 1, 99, 2, 
/* out0334_em-eta2-phi8 */     1, 35, 1, 
/* out0335_em-eta2-phi9 */     2, 35, 3, 37, 1, 
/* out0336_em-eta1-phi10 */     2, 37, 1, 72, 4, 
/* out0337_em-eta1-phi11 */     1, 72, 2, 
/* out0338_em-eta0-phi12 */     0, 
/* out0339_em-eta0-phi13 */     2, 62, 2, 105, 1, 
/* out0340_em-eta0-phi0 */     1, 36, 3, 
/* out0341_em-eta0-phi1 */     0, 
/* out0342_em-eta0-phi2 */     2, 7, 1, 48, 1, 
/* out0343_em-eta1-phi2 */     3, 7, 5, 48, 1, 80, 1, 
/* out0344_em-eta1-phi3 */     4, 7, 1, 47, 2, 48, 3, 80, 6, 
/* out0345_em-eta1-phi4 */     1, 47, 1, 
/* out0346_em-eta1-phi5 */     1, 21, 2, 
/* out0347_em-eta1-phi6 */     5, 20, 3, 21, 2, 22, 1, 64, 2, 99, 1, 
/* out0348_em-eta1-phi7 */     5, 20, 1, 22, 2, 64, 5, 99, 5, 100, 1, 
/* out0349_em-eta1-phi8 */     1, 37, 1, 
/* out0350_em-eta0-phi9 */     1, 38, 5, 
/* out0351_em-eta1-phi9 */     1, 37, 5, 
/* out0352_em-eta0-phi10 */     1, 38, 3, 
/* out0353_em-eta0-phi11 */     0, 
/* out0354_em-eta0-phi3 */     2, 48, 3, 80, 1, 
/* out0355_em-eta0-phi4 */     0, 
/* out0356_em-eta0-phi5 */     1, 21, 2, 
/* out0357_em-eta0-phi6 */     2, 21, 2, 22, 1, 
/* out0358_em-eta0-phi7 */     3, 22, 4, 64, 1, 100, 5, 
/* out0359_em-eta0-phi8 */     1, 100, 2, 
/* out0360_em-eta17-phi19 */     0, 
/* out0361_em-eta17-phi20 */     0, 
/* out0362_em-eta16-phi-2 */     0, 
/* out0363_em-eta16-phi1 */     0, 
/* out0364_em-eta17-phi0 */     0, 
/* out0365_em-eta17-phi3 */     1, 13, 1, 
/* out0366_em-eta17-phi4 */     2, 13, 1, 65, 1, 
/* out0367_em-eta16-phi11 */     1, 66, 1, 
/* out0368_em-eta14-phi14 */     1, 8, 1, 
/* out0369_em-eta14-phi15 */     0, 
/* out0370_em-eta11-phi16 */     1, 49, 1, 
/* out0371_em-eta13-phi-1 */     0, 
/* out0372_em-eta14-phi8 */     1, 67, 1, 
/* out0373_em-eta14-phi9 */     1, 67, 1, 
/* out0374_em-eta9-phi-2 */     0, 
/* out0375_em-eta11-phi7 */     1, 39, 1, 
/* out0376_em-eta14-phi19 */     1, 82, 1, 
/* out0377_em-eta14-phi17 */     1, 8, 1, 
/* out0378_em-eta11-phi19 */     1, 49, 1, 
/* out0379_em-eta14-phi4 */     2, 14, 1, 42, 1, 
/* out0380_em-eta14-phi6 */     1, 67, 1, 
/* out0381_em-eta11-phi4 */     1, 39, 1, 
/* out0382_em-eta14-phi21 */     1, 82, 1, 
/* out0383_em-eta11-phi22 */     1, 83, 1, 
/* out0384_em-eta12-phi17 */     1, 49, 1, 
/* out0385_em-eta14-phi2 */     2, 14, 1, 42, 1, 
/* out0386_em-eta11-phi13 */     0, 
/* out0387_em-eta12-phi6 */     1, 39, 1, 
/* out0388_em-eta11-phi10 */     0, 
/* out0389_em-eta4-phi23 */     2, 74, 1, 85, 1, 
/* out0390_em-eta17-phi11 */     1, 66, 1, 
/* out0391_em-eta12-phi18 */     1, 49, 1, 
/* out0392_em-eta12-phi5 */     1, 39, 1, 
/* out0393_em-eta0-phi-1 */     1, 36, 3, 
/* out0394_em-eta14-phi18 */     1, 82, 1, 
/* out0395_em-eta6-phi23 */     2, 73, 1, 84, 1, 
/* out0396_em-eta17-phi13 */     1, 66, 1, 
/* out0397_em-eta14-phi5 */     1, 42, 1, 
/* out0398_em-eta17-phi2 */     0, 
/* out0399_em-eta17-phi-2 */     0, 
/* out0400_em-eta17-phi1 */     0, 
/* out0401_em-eta17-phi10 */     1, 66, 1, 
/* out0402_em-eta15-phi15 */     0, 
/* out0403_em-eta14-phi0 */     0, 
/* out0404_em-eta15-phi8 */     0, 
/* out0405_em-eta13-phi10 */     1, 68, 1, 
/* out0406_em-eta13-phi13 */     1, 68, 1, 
/* out0407_em-eta15-phi20 */     0, 
/* out0408_em-eta17-phi-3 */     0, 
/* out0409_em-eta17-phi-1 */     0, 
/* out0410_em-eta15-phi16 */     0, 
/* out0411_em-eta13-phi-2 */     0, 
/* out0412_em-eta13-phi1 */     0, 
/* out0413_em-eta15-phi3 */     0, 
/* out0414_em-eta15-phi7 */     1, 67, 1, 
/* out0415_em-eta14-phi11 */     0, 
/* out0416_em-eta14-phi12 */     1, 68, 1, 
/* out0417_em-eta14-phi-1 */     0, 
/* out0418_em-eta15-phi14 */     0, 
/* out0419_em-eta15-phi9 */     0, 
/* out0420_em-eta10-phi-2 */     0, 
/* out0421_em-eta15-phi19 */     1, 82, 1, 
/* out0422_em-eta15-phi21 */     1, 82, 1, 
/* out0423_em-eta15-phi17 */     0, 
/* out0424_em-eta15-phi2 */     0, 
/* out0425_em-eta15-phi4 */     0, 
/* out0426_em-eta15-phi6 */     0, 
/* out0427_em-eta12-phi22 */     0
};