parameter integer matrixE [0:1587] = {
/* num inputs = 117 (in0-in116) */
/* num outputs = 428(out0-out427) */
//* max inputs per outputs = 6 */
//* total number of input in adders 580 */

/* out0000_em-eta16-phi16 */     0, 
/* out0001_em-eta16-phi17 */     2, 11, 1, 46, 1, 
/* out0002_em-eta16-phi18 */     1, 11, 1, 
/* out0003_em-eta16-phi19 */     0, 
/* out0004_em-eta17-phi15 */     0, 
/* out0005_em-eta17-phi16 */     2, 11, 1, 46, 1, 
/* out0006_em-eta17-phi17 */     2, 11, 1, 46, 1, 
/* out0007_em-eta17-phi18 */     2, 11, 1, 46, 1, 
/* out0008_em-eta12-phi19 */     2, 26, 1, 103, 1, 
/* out0009_em-eta12-phi20 */     0, 
/* out0010_em-eta12-phi21 */     1, 48, 1, 
/* out0011_em-eta13-phi18 */     2, 26, 1, 47, 1, 
/* out0012_em-eta13-phi19 */     2, 26, 1, 47, 1, 
/* out0013_em-eta13-phi20 */     2, 26, 1, 47, 1, 
/* out0014_em-eta13-phi21 */     2, 26, 1, 47, 1, 
/* out0015_em-eta14-phi20 */     2, 26, 1, 47, 1, 
/* out0016_em-eta9-phi20 */     3, 27, 1, 30, 1, 104, 1, 
/* out0017_em-eta9-phi21 */     3, 27, 1, 48, 1, 49, 1, 
/* out0018_em-eta9-phi22 */     1, 49, 1, 
/* out0019_em-eta10-phi20 */     2, 27, 1, 48, 1, 
/* out0020_em-eta10-phi21 */     2, 27, 1, 48, 1, 
/* out0021_em-eta10-phi22 */     2, 27, 1, 48, 1, 
/* out0022_em-eta11-phi20 */     2, 27, 1, 48, 1, 
/* out0023_em-eta11-phi21 */     2, 27, 1, 48, 1, 
/* out0024_em-eta6-phi21 */     1, 0, 1, 
/* out0025_em-eta6-phi22 */     2, 0, 1, 1, 1, 
/* out0026_em-eta7-phi20 */     1, 0, 1, 
/* out0027_em-eta7-phi21 */     2, 0, 1, 49, 1, 
/* out0028_em-eta7-phi22 */     2, 0, 2, 49, 1, 
/* out0029_em-eta8-phi21 */     2, 0, 1, 49, 2, 
/* out0030_em-eta8-phi22 */     2, 0, 1, 49, 1, 
/* out0031_em-eta4-phi21 */     1, 1, 1, 
/* out0032_em-eta4-phi22 */     1, 1, 1, 
/* out0033_em-eta5-phi21 */     1, 1, 2, 
/* out0034_em-eta5-phi22 */     1, 1, 2, 
/* out0035_em-eta5-phi23 */     1, 1, 1, 
/* out0036_em-eta2-phi22 */     0, 
/* out0037_em-eta3-phi21 */     0, 
/* out0038_em-eta3-phi22 */     0, 
/* out0039_em-eta3-phi23 */     0, 
/* out0040_em-eta1-phi22 */     1, 19, 3, 
/* out0041_em-eta1-phi23 */     1, 19, 2, 
/* out0042_em-eta2-phi23 */     0, 
/* out0043_em-eta0-phi22 */     1, 19, 2, 
/* out0044_em-eta0-phi23 */     1, 19, 1, 
/* out0045_em-eta15-phi-2 */     1, 20, 1, 
/* out0046_em-eta15-phi-1 */     1, 20, 1, 
/* out0047_em-eta15-phi0 */     1, 20, 1, 
/* out0048_em-eta15-phi1 */     1, 20, 1, 
/* out0049_em-eta16-phi-3 */     0, 
/* out0050_em-eta16-phi-1 */     0, 
/* out0051_em-eta16-phi0 */     1, 20, 1, 
/* out0052_em-eta16-phi2 */     0, 
/* out0053_em-eta16-phi4 */     0, 
/* out0054_em-eta16-phi5 */     0, 
/* out0055_em-eta16-phi6 */     0, 
/* out0056_em-eta16-phi7 */     0, 
/* out0057_em-eta17-phi5 */     1, 102, 1, 
/* out0058_em-eta17-phi6 */     1, 102, 1, 
/* out0059_em-eta17-phi7 */     0, 
/* out0060_em-eta17-phi8 */     0, 
/* out0061_em-eta15-phi10 */     0, 
/* out0062_em-eta15-phi11 */     0, 
/* out0063_em-eta15-phi12 */     0, 
/* out0064_em-eta15-phi13 */     0, 
/* out0065_em-eta16-phi10 */     0, 
/* out0066_em-eta16-phi12 */     0, 
/* out0067_em-eta16-phi13 */     0, 
/* out0068_em-eta17-phi12 */     0, 
/* out0069_em-eta12-phi14 */     0, 
/* out0070_em-eta12-phi15 */     0, 
/* out0071_em-eta12-phi16 */     1, 103, 1, 
/* out0072_em-eta13-phi14 */     0, 
/* out0073_em-eta13-phi15 */     0, 
/* out0074_em-eta13-phi16 */     0, 
/* out0075_em-eta13-phi17 */     0, 
/* out0076_em-eta14-phi16 */     0, 
/* out0077_em-eta9-phi17 */     2, 31, 1, 106, 1, 
/* out0078_em-eta9-phi18 */     2, 30, 1, 104, 1, 
/* out0079_em-eta10-phi16 */     1, 106, 1, 
/* out0080_em-eta10-phi17 */     3, 29, 1, 103, 1, 106, 1, 
/* out0081_em-eta10-phi18 */     2, 29, 1, 104, 1, 
/* out0082_em-eta10-phi19 */     1, 104, 1, 
/* out0083_em-eta11-phi17 */     2, 29, 1, 103, 1, 
/* out0084_em-eta11-phi18 */     2, 29, 1, 103, 1, 
/* out0085_em-eta7-phi18 */     1, 32, 1, 
/* out0086_em-eta7-phi19 */     1, 30, 1, 
/* out0087_em-eta8-phi18 */     2, 30, 1, 104, 1, 
/* out0088_em-eta8-phi19 */     2, 30, 2, 104, 1, 
/* out0089_em-eta8-phi20 */     3, 30, 1, 49, 1, 104, 1, 
/* out0090_em-eta9-phi19 */     2, 30, 1, 104, 1, 
/* out0091_em-eta5-phi19 */     1, 33, 2, 
/* out0092_em-eta5-phi20 */     0, 
/* out0093_em-eta6-phi19 */     0, 
/* out0094_em-eta6-phi20 */     0, 
/* out0095_em-eta3-phi20 */     1, 34, 2, 
/* out0096_em-eta4-phi20 */     0, 
/* out0097_em-eta2-phi20 */     0, 
/* out0098_em-eta2-phi21 */     0, 
/* out0099_em-eta0-phi21 */     0, 
/* out0100_em-eta1-phi21 */     0, 
/* out0101_em-eta11-phi-1 */     2, 21, 1, 75, 1, 
/* out0102_em-eta11-phi0 */     2, 21, 1, 75, 1, 
/* out0103_em-eta11-phi1 */     0, 
/* out0104_em-eta12-phi-2 */     1, 21, 1, 
/* out0105_em-eta12-phi-1 */     1, 21, 1, 
/* out0106_em-eta12-phi0 */     1, 21, 1, 
/* out0107_em-eta12-phi1 */     1, 21, 1, 
/* out0108_em-eta13-phi0 */     1, 21, 1, 
/* out0109_em-eta12-phi2 */     0, 
/* out0110_em-eta12-phi3 */     0, 
/* out0111_em-eta12-phi4 */     1, 109, 1, 
/* out0112_em-eta13-phi2 */     0, 
/* out0113_em-eta13-phi3 */     0, 
/* out0114_em-eta13-phi4 */     0, 
/* out0115_em-eta13-phi5 */     0, 
/* out0116_em-eta14-phi3 */     0, 
/* out0117_em-eta12-phi7 */     1, 109, 1, 
/* out0118_em-eta12-phi8 */     2, 76, 1, 107, 1, 
/* out0119_em-eta12-phi9 */     2, 76, 1, 107, 1, 
/* out0120_em-eta13-phi6 */     1, 109, 1, 
/* out0121_em-eta13-phi7 */     1, 105, 1, 
/* out0122_em-eta13-phi8 */     1, 105, 1, 
/* out0123_em-eta13-phi9 */     0, 
/* out0124_em-eta14-phi7 */     1, 105, 1, 
/* out0125_em-eta11-phi11 */     0, 
/* out0126_em-eta11-phi12 */     0, 
/* out0127_em-eta12-phi10 */     0, 
/* out0128_em-eta12-phi11 */     0, 
/* out0129_em-eta12-phi12 */     0, 
/* out0130_em-eta12-phi13 */     0, 
/* out0131_em-eta13-phi11 */     0, 
/* out0132_em-eta13-phi12 */     0, 
/* out0133_em-eta9-phi13 */     0, 
/* out0134_em-eta9-phi14 */     0, 
/* out0135_em-eta9-phi15 */     2, 31, 1, 106, 1, 
/* out0136_em-eta10-phi13 */     0, 
/* out0137_em-eta10-phi14 */     0, 
/* out0138_em-eta10-phi15 */     0, 
/* out0139_em-eta11-phi14 */     0, 
/* out0140_em-eta11-phi15 */     0, 
/* out0141_em-eta7-phi15 */     1, 12, 1, 
/* out0142_em-eta7-phi16 */     1, 31, 1, 
/* out0143_em-eta7-phi17 */     1, 32, 2, 
/* out0144_em-eta8-phi15 */     2, 31, 1, 106, 1, 
/* out0145_em-eta8-phi16 */     2, 31, 2, 106, 1, 
/* out0146_em-eta8-phi17 */     2, 31, 1, 106, 1, 
/* out0147_em-eta9-phi16 */     2, 31, 1, 106, 1, 
/* out0148_em-eta5-phi17 */     1, 32, 1, 
/* out0149_em-eta5-phi18 */     1, 33, 2, 
/* out0150_em-eta6-phi17 */     1, 32, 2, 
/* out0151_em-eta6-phi18 */     1, 32, 2, 
/* out0152_em-eta3-phi18 */     5, 13, 3, 50, 3, 51, 1, 77, 2, 78, 1, 
/* out0153_em-eta3-phi19 */     2, 34, 4, 78, 1, 
/* out0154_em-eta4-phi18 */     3, 33, 2, 50, 1, 77, 2, 
/* out0155_em-eta4-phi19 */     2, 33, 2, 34, 1, 
/* out0156_em-eta2-phi19 */     4, 34, 1, 51, 2, 78, 2, 79, 1, 
/* out0157_em-eta1-phi19 */     2, 52, 5, 79, 5, 
/* out0158_em-eta1-phi20 */     0, 
/* out0159_em-eta0-phi20 */     0, 
/* out0160_em-eta8-phi-1 */     2, 22, 1, 53, 1, 
/* out0161_em-eta8-phi0 */     2, 22, 1, 53, 1, 
/* out0162_em-eta9-phi-1 */     2, 22, 1, 75, 1, 
/* out0163_em-eta9-phi0 */     2, 22, 1, 75, 2, 
/* out0164_em-eta9-phi1 */     1, 22, 1, 
/* out0165_em-eta10-phi-1 */     2, 22, 1, 75, 1, 
/* out0166_em-eta10-phi0 */     2, 22, 1, 75, 1, 
/* out0167_em-eta9-phi2 */     0, 
/* out0168_em-eta9-phi3 */     1, 110, 1, 
/* out0169_em-eta10-phi1 */     1, 75, 1, 
/* out0170_em-eta10-phi2 */     0, 
/* out0171_em-eta10-phi3 */     0, 
/* out0172_em-eta11-phi2 */     0, 
/* out0173_em-eta11-phi3 */     0, 
/* out0174_em-eta9-phi5 */     1, 110, 1, 
/* out0175_em-eta9-phi6 */     2, 45, 1, 111, 1, 
/* out0176_em-eta10-phi4 */     1, 110, 1, 
/* out0177_em-eta10-phi5 */     2, 44, 1, 110, 1, 
/* out0178_em-eta10-phi6 */     2, 44, 1, 111, 1, 
/* out0179_em-eta10-phi7 */     1, 111, 1, 
/* out0180_em-eta11-phi5 */     2, 44, 1, 109, 1, 
/* out0181_em-eta11-phi6 */     2, 44, 1, 109, 1, 
/* out0182_em-eta9-phi8 */     2, 45, 1, 111, 1, 
/* out0183_em-eta9-phi9 */     3, 80, 1, 91, 1, 108, 1, 
/* out0184_em-eta9-phi10 */     3, 80, 1, 91, 1, 108, 1, 
/* out0185_em-eta10-phi8 */     2, 76, 1, 107, 1, 
/* out0186_em-eta10-phi9 */     2, 76, 1, 107, 1, 
/* out0187_em-eta10-phi10 */     2, 76, 1, 107, 1, 
/* out0188_em-eta11-phi8 */     2, 76, 1, 107, 1, 
/* out0189_em-eta11-phi9 */     2, 76, 1, 107, 1, 
/* out0190_em-eta8-phi11 */     1, 54, 1, 
/* out0191_em-eta8-phi12 */     1, 54, 1, 
/* out0192_em-eta9-phi11 */     0, 
/* out0193_em-eta9-phi12 */     0, 
/* out0194_em-eta10-phi11 */     0, 
/* out0195_em-eta10-phi12 */     0, 
/* out0196_em-eta6-phi13 */     1, 81, 2, 
/* out0197_em-eta6-phi14 */     1, 81, 2, 
/* out0198_em-eta7-phi13 */     1, 81, 1, 
/* out0199_em-eta7-phi14 */     0, 
/* out0200_em-eta8-phi13 */     0, 
/* out0201_em-eta8-phi14 */     0, 
/* out0202_em-eta5-phi15 */     2, 12, 2, 14, 1, 
/* out0203_em-eta5-phi16 */     1, 12, 1, 
/* out0204_em-eta6-phi15 */     1, 12, 2, 
/* out0205_em-eta6-phi16 */     1, 12, 2, 
/* out0206_em-eta3-phi16 */     0, 
/* out0207_em-eta3-phi17 */     3, 13, 3, 50, 3, 77, 2, 
/* out0208_em-eta4-phi16 */     0, 
/* out0209_em-eta4-phi17 */     2, 50, 1, 77, 2, 
/* out0210_em-eta2-phi17 */     2, 13, 1, 15, 3, 
/* out0211_em-eta2-phi18 */     3, 13, 1, 51, 4, 78, 4, 
/* out0212_em-eta1-phi18 */     3, 51, 1, 52, 1, 79, 2, 
/* out0213_em-eta0-phi18 */     0, 
/* out0214_em-eta0-phi19 */     1, 52, 2, 
/* out0215_em-eta5-phi-1 */     2, 36, 2, 55, 2, 
/* out0216_em-eta5-phi0 */     2, 36, 2, 55, 3, 
/* out0217_em-eta6-phi-1 */     2, 35, 2, 53, 1, 
/* out0218_em-eta6-phi0 */     5, 35, 2, 37, 1, 53, 1, 55, 1, 82, 1, 
/* out0219_em-eta7-phi-1 */     2, 35, 2, 53, 2, 
/* out0220_em-eta7-phi0 */     2, 35, 2, 53, 2, 
/* out0221_em-eta6-phi1 */     2, 37, 2, 82, 2, 
/* out0222_em-eta6-phi2 */     2, 37, 1, 82, 2, 
/* out0223_em-eta7-phi1 */     1, 82, 1, 
/* out0224_em-eta7-phi2 */     1, 112, 1, 
/* out0225_em-eta7-phi3 */     2, 92, 2, 112, 2, 
/* out0226_em-eta8-phi1 */     0, 
/* out0227_em-eta8-phi2 */     0, 
/* out0228_em-eta7-phi4 */     2, 92, 2, 112, 2, 
/* out0229_em-eta7-phi5 */     2, 67, 2, 93, 2, 
/* out0230_em-eta8-phi3 */     2, 110, 1, 112, 1, 
/* out0231_em-eta8-phi4 */     1, 110, 1, 
/* out0232_em-eta8-phi5 */     1, 110, 1, 
/* out0233_em-eta9-phi4 */     1, 110, 1, 
/* out0234_em-eta7-phi6 */     3, 3, 1, 67, 2, 93, 2, 
/* out0235_em-eta7-phi7 */     1, 45, 1, 
/* out0236_em-eta7-phi8 */     0, 
/* out0237_em-eta8-phi6 */     3, 45, 1, 93, 1, 111, 1, 
/* out0238_em-eta8-phi7 */     2, 45, 2, 111, 1, 
/* out0239_em-eta8-phi8 */     4, 45, 1, 80, 1, 91, 1, 108, 1, 
/* out0240_em-eta9-phi7 */     2, 45, 1, 111, 2, 
/* out0241_em-eta6-phi9 */     0, 
/* out0242_em-eta6-phi10 */     0, 
/* out0243_em-eta7-phi9 */     3, 80, 1, 91, 1, 108, 1, 
/* out0244_em-eta7-phi10 */     2, 80, 1, 91, 1, 
/* out0245_em-eta8-phi9 */     3, 80, 2, 91, 2, 108, 2, 
/* out0246_em-eta8-phi10 */     3, 80, 1, 91, 1, 108, 2, 
/* out0247_em-eta5-phi11 */     3, 2, 1, 4, 1, 56, 2, 
/* out0248_em-eta5-phi12 */     3, 2, 1, 4, 1, 56, 3, 
/* out0249_em-eta6-phi11 */     2, 2, 2, 54, 1, 
/* out0250_em-eta6-phi12 */     4, 2, 2, 54, 1, 56, 1, 81, 1, 
/* out0251_em-eta7-phi11 */     2, 2, 1, 54, 2, 
/* out0252_em-eta7-phi12 */     2, 2, 1, 54, 2, 
/* out0253_em-eta4-phi13 */     1, 83, 3, 
/* out0254_em-eta4-phi14 */     2, 14, 2, 83, 1, 
/* out0255_em-eta5-phi13 */     2, 81, 1, 83, 2, 
/* out0256_em-eta5-phi14 */     1, 81, 1, 
/* out0257_em-eta3-phi14 */     2, 14, 1, 16, 2, 
/* out0258_em-eta3-phi15 */     2, 14, 1, 16, 1, 
/* out0259_em-eta4-phi15 */     1, 14, 3, 
/* out0260_em-eta2-phi15 */     1, 16, 2, 
/* out0261_em-eta2-phi16 */     1, 15, 1, 
/* out0262_em-eta1-phi16 */     2, 15, 1, 17, 2, 
/* out0263_em-eta1-phi17 */     2, 15, 3, 17, 1, 
/* out0264_em-eta0-phi17 */     1, 17, 1, 
/* out0265_em-eta3-phi0 */     3, 38, 3, 57, 3, 86, 1, 
/* out0266_em-eta4-phi-1 */     3, 36, 2, 55, 1, 57, 1, 
/* out0267_em-eta4-phi0 */     5, 36, 2, 39, 1, 55, 1, 57, 1, 84, 1, 
/* out0268_em-eta4-phi1 */     2, 39, 3, 84, 3, 
/* out0269_em-eta4-phi2 */     6, 39, 1, 84, 1, 94, 1, 96, 1, 113, 1, 114, 2, 
/* out0270_em-eta5-phi1 */     3, 37, 2, 82, 1, 84, 2, 
/* out0271_em-eta5-phi2 */     4, 37, 2, 82, 1, 94, 2, 113, 2, 
/* out0272_em-eta5-phi3 */     2, 94, 3, 113, 3, 
/* out0273_em-eta5-phi4 */     1, 58, 2, 
/* out0274_em-eta6-phi3 */     3, 92, 2, 112, 1, 113, 1, 
/* out0275_em-eta6-phi4 */     2, 92, 2, 112, 1, 
/* out0276_em-eta5-phi5 */     2, 3, 1, 58, 2, 
/* out0277_em-eta5-phi6 */     4, 3, 2, 5, 1, 68, 3, 95, 3, 
/* out0278_em-eta6-phi5 */     3, 3, 2, 67, 2, 93, 1, 
/* out0279_em-eta6-phi6 */     4, 3, 2, 67, 2, 93, 2, 95, 1, 
/* out0280_em-eta5-phi7 */     2, 68, 2, 95, 2, 
/* out0281_em-eta5-phi8 */     0, 
/* out0282_em-eta6-phi7 */     1, 95, 1, 
/* out0283_em-eta6-phi8 */     0, 
/* out0284_em-eta4-phi9 */     0, 
/* out0285_em-eta4-phi10 */     0, 
/* out0286_em-eta5-phi9 */     0, 
/* out0287_em-eta5-phi10 */     0, 
/* out0288_em-eta3-phi12 */     4, 4, 1, 6, 2, 59, 3, 85, 1, 
/* out0289_em-eta4-phi11 */     3, 4, 2, 56, 1, 59, 1, 
/* out0290_em-eta4-phi12 */     4, 4, 3, 56, 1, 59, 1, 83, 1, 
/* out0291_em-eta2-phi13 */     2, 85, 3, 87, 1, 
/* out0292_em-eta3-phi13 */     2, 83, 1, 85, 3, 
/* out0293_em-eta2-phi14 */     1, 16, 3, 
/* out0294_em-eta1-phi15 */     2, 18, 1, 28, 2, 
/* out0295_em-eta0-phi16 */     1, 17, 4, 
/* out0296_em-eta2-phi-1 */     3, 38, 1, 40, 2, 60, 2, 
/* out0297_em-eta2-phi0 */     6, 38, 1, 40, 2, 41, 2, 60, 3, 86, 1, 88, 1, 
/* out0298_em-eta3-phi-1 */     2, 38, 3, 57, 3, 
/* out0299_em-eta2-phi1 */     5, 41, 4, 86, 3, 88, 1, 98, 1, 115, 1, 
/* out0300_em-eta3-phi1 */     4, 39, 2, 41, 1, 84, 1, 86, 3, 
/* out0301_em-eta3-phi2 */     4, 39, 1, 96, 4, 114, 3, 115, 1, 
/* out0302_em-eta3-phi3 */     3, 61, 2, 96, 2, 114, 2, 
/* out0303_em-eta4-phi3 */     4, 94, 2, 96, 1, 113, 1, 114, 1, 
/* out0304_em-eta3-phi4 */     1, 61, 4, 
/* out0305_em-eta3-phi5 */     3, 23, 3, 61, 1, 72, 1, 
/* out0306_em-eta4-phi4 */     2, 58, 2, 61, 1, 
/* out0307_em-eta4-phi5 */     1, 58, 2, 
/* out0308_em-eta3-phi6 */     2, 5, 1, 23, 3, 
/* out0309_em-eta3-phi7 */     5, 5, 1, 7, 3, 69, 4, 97, 3, 99, 1, 
/* out0310_em-eta4-phi6 */     3, 5, 3, 68, 2, 95, 1, 
/* out0311_em-eta4-phi7 */     4, 5, 2, 68, 1, 69, 2, 97, 3, 
/* out0312_em-eta3-phi8 */     4, 7, 1, 69, 1, 97, 1, 99, 1, 
/* out0313_em-eta3-phi9 */     0, 
/* out0314_em-eta4-phi8 */     2, 69, 1, 97, 1, 
/* out0315_em-eta2-phi10 */     0, 
/* out0316_em-eta3-phi10 */     0, 
/* out0317_em-eta3-phi11 */     2, 6, 2, 59, 3, 
/* out0318_em-eta2-phi11 */     2, 6, 2, 62, 3, 
/* out0319_em-eta2-phi12 */     5, 6, 2, 8, 1, 62, 3, 85, 1, 87, 1, 
/* out0320_em-eta1-phi12 */     4, 8, 3, 62, 1, 65, 2, 87, 2, 
/* out0321_em-eta1-phi13 */     3, 18, 1, 87, 4, 89, 1, 
/* out0322_em-eta0-phi14 */     2, 18, 1, 28, 1, 
/* out0323_em-eta1-phi14 */     1, 18, 5, 
/* out0324_em-eta0-phi15 */     1, 28, 5, 
/* out0325_em-eta1-phi-1 */     4, 40, 2, 42, 1, 60, 1, 63, 2, 
/* out0326_em-eta1-phi0 */     6, 40, 2, 42, 1, 43, 2, 60, 2, 63, 2, 88, 2, 
/* out0327_em-eta1-phi1 */     5, 43, 4, 88, 4, 90, 1, 100, 2, 116, 2, 
/* out0328_em-eta2-phi2 */     3, 41, 1, 98, 5, 115, 5, 
/* out0329_em-eta2-phi3 */     1, 64, 4, 
/* out0330_em-eta2-phi4 */     3, 24, 1, 64, 2, 72, 2, 
/* out0331_em-eta2-phi5 */     3, 23, 1, 24, 3, 72, 5, 
/* out0332_em-eta2-phi6 */     1, 23, 1, 
/* out0333_em-eta2-phi7 */     3, 7, 3, 70, 2, 99, 2, 
/* out0334_em-eta2-phi8 */     4, 7, 1, 9, 1, 70, 4, 99, 4, 
/* out0335_em-eta2-phi9 */     0, 
/* out0336_em-eta1-phi10 */     0, 
/* out0337_em-eta1-phi11 */     3, 8, 3, 62, 1, 65, 2, 
/* out0338_em-eta0-phi12 */     3, 8, 1, 65, 2, 89, 3, 
/* out0339_em-eta0-phi13 */     1, 89, 4, 
/* out0340_em-eta0-phi0 */     4, 42, 3, 43, 1, 63, 2, 90, 3, 
/* out0341_em-eta0-phi1 */     4, 43, 1, 90, 4, 100, 1, 116, 1, 
/* out0342_em-eta0-phi2 */     2, 100, 2, 116, 1, 
/* out0343_em-eta1-phi2 */     5, 66, 1, 98, 2, 100, 3, 115, 1, 116, 4, 
/* out0344_em-eta1-phi3 */     2, 64, 1, 66, 4, 
/* out0345_em-eta1-phi4 */     4, 24, 1, 25, 2, 64, 1, 73, 5, 
/* out0346_em-eta1-phi5 */     4, 24, 3, 25, 1, 73, 2, 74, 4, 
/* out0347_em-eta1-phi6 */     1, 74, 4, 
/* out0348_em-eta1-phi7 */     2, 9, 3, 70, 1, 
/* out0349_em-eta1-phi8 */     4, 9, 4, 70, 1, 71, 4, 101, 6, 
/* out0350_em-eta0-phi9 */     1, 10, 1, 
/* out0351_em-eta1-phi9 */     2, 71, 1, 101, 1, 
/* out0352_em-eta0-phi10 */     0, 
/* out0353_em-eta0-phi11 */     1, 65, 2, 
/* out0354_em-eta0-phi3 */     1, 66, 3, 
/* out0355_em-eta0-phi4 */     2, 25, 4, 73, 1, 
/* out0356_em-eta0-phi5 */     1, 25, 1, 
/* out0357_em-eta0-phi6 */     0, 
/* out0358_em-eta0-phi7 */     0, 
/* out0359_em-eta0-phi8 */     3, 10, 7, 71, 3, 101, 1, 
/* out0360_em-eta17-phi19 */     2, 11, 1, 46, 1, 
/* out0361_em-eta17-phi20 */     1, 11, 1, 
/* out0362_em-eta16-phi-2 */     1, 20, 1, 
/* out0363_em-eta16-phi1 */     1, 20, 1, 
/* out0364_em-eta17-phi0 */     1, 20, 1, 
/* out0365_em-eta17-phi3 */     0, 
/* out0366_em-eta17-phi4 */     0, 
/* out0367_em-eta16-phi11 */     0, 
/* out0368_em-eta14-phi14 */     0, 
/* out0369_em-eta14-phi15 */     0, 
/* out0370_em-eta11-phi16 */     1, 29, 1, 
/* out0371_em-eta13-phi-1 */     1, 21, 1, 
/* out0372_em-eta14-phi8 */     1, 105, 1, 
/* out0373_em-eta14-phi9 */     1, 105, 1, 
/* out0374_em-eta9-phi-2 */     1, 22, 1, 
/* out0375_em-eta11-phi7 */     1, 44, 1, 
/* out0376_em-eta14-phi19 */     2, 26, 1, 47, 1, 
/* out0377_em-eta14-phi17 */     0, 
/* out0378_em-eta11-phi19 */     2, 29, 1, 103, 1, 
/* out0379_em-eta14-phi4 */     0, 
/* out0380_em-eta14-phi6 */     1, 105, 1, 
/* out0381_em-eta11-phi4 */     2, 44, 1, 109, 1, 
/* out0382_em-eta14-phi21 */     2, 26, 1, 47, 1, 
/* out0383_em-eta11-phi22 */     2, 27, 1, 48, 1, 
/* out0384_em-eta12-phi17 */     2, 29, 1, 103, 1, 
/* out0385_em-eta14-phi2 */     0, 
/* out0386_em-eta11-phi13 */     0, 
/* out0387_em-eta12-phi6 */     2, 44, 1, 109, 1, 
/* out0388_em-eta11-phi10 */     2, 76, 1, 107, 1, 
/* out0389_em-eta4-phi23 */     0, 
/* out0390_em-eta17-phi11 */     0, 
/* out0391_em-eta12-phi18 */     2, 29, 1, 103, 1, 
/* out0392_em-eta12-phi5 */     2, 44, 1, 109, 1, 
/* out0393_em-eta0-phi-1 */     2, 42, 3, 63, 2, 
/* out0394_em-eta14-phi18 */     1, 47, 1, 
/* out0395_em-eta6-phi23 */     0, 
/* out0396_em-eta17-phi13 */     0, 
/* out0397_em-eta14-phi5 */     0, 
/* out0398_em-eta17-phi2 */     0, 
/* out0399_em-eta17-phi-2 */     0, 
/* out0400_em-eta17-phi1 */     0, 
/* out0401_em-eta17-phi10 */     0, 
/* out0402_em-eta15-phi15 */     0, 
/* out0403_em-eta14-phi0 */     0, 
/* out0404_em-eta15-phi8 */     0, 
/* out0405_em-eta13-phi10 */     0, 
/* out0406_em-eta13-phi13 */     0, 
/* out0407_em-eta15-phi20 */     0, 
/* out0408_em-eta17-phi-3 */     0, 
/* out0409_em-eta17-phi-1 */     0, 
/* out0410_em-eta15-phi16 */     0, 
/* out0411_em-eta13-phi-2 */     0, 
/* out0412_em-eta13-phi1 */     0, 
/* out0413_em-eta15-phi3 */     0, 
/* out0414_em-eta15-phi7 */     0, 
/* out0415_em-eta14-phi11 */     0, 
/* out0416_em-eta14-phi12 */     0, 
/* out0417_em-eta14-phi-1 */     0, 
/* out0418_em-eta15-phi14 */     0, 
/* out0419_em-eta15-phi9 */     1, 105, 1, 
/* out0420_em-eta10-phi-2 */     0, 
/* out0421_em-eta15-phi19 */     0, 
/* out0422_em-eta15-phi21 */     0, 
/* out0423_em-eta15-phi17 */     0, 
/* out0424_em-eta15-phi2 */     0, 
/* out0425_em-eta15-phi4 */     0, 
/* out0426_em-eta15-phi6 */     1, 105, 1, 
/* out0427_em-eta12-phi22 */     0
};