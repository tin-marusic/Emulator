parameter integer matrixH [0:2454] = {
/* num inputs = 192 (in0-in191) */
/* num outputs = 515(out0-out514) */
//* max inputs per outputs = 14 */
//* total number of input in adders 970 */

/* out0000_had-eta14-phi21 */     4, 114, 2, 119, 2, 138, 2, 159, 2, 
/* out0001_had-eta14-phi22 */     4, 119, 2, 134, 2, 148, 2, 159, 2, 
/* out0002_had-eta14-phi23 */     4, 119, 2, 134, 2, 148, 2, 159, 2, 
/* out0003_had-eta15-phi21 */     4, 114, 2, 134, 2, 148, 2, 159, 2, 
/* out0004_had-eta15-phi22 */     4, 119, 2, 134, 2, 148, 2, 159, 2, 
/* out0005_had-eta15-phi23 */     3, 119, 2, 134, 2, 148, 2, 
/* out0006_had-eta15-phi24 */     2, 134, 2, 148, 2, 
/* out0007_had-eta16-phi22 */     3, 134, 2, 148, 2, 158, 2, 
/* out0008_had-eta11-phi22 */     5, 120, 2, 135, 2, 139, 2, 150, 2, 160, 4, 
/* out0009_had-eta11-phi23 */     6, 120, 4, 135, 2, 136, 2, 149, 2, 150, 2, 160, 2, 
/* out0010_had-eta11-phi24 */     0, 
/* out0011_had-eta12-phi22 */     4, 120, 2, 135, 4, 149, 4, 160, 4, 
/* out0012_had-eta12-phi23 */     4, 120, 4, 135, 2, 149, 4, 160, 2, 
/* out0013_had-eta12-phi24 */     3, 120, 2, 135, 2, 149, 2, 
/* out0014_had-eta13-phi22 */     4, 119, 2, 135, 2, 149, 2, 159, 2, 
/* out0015_had-eta13-phi23 */     5, 119, 2, 120, 2, 135, 2, 149, 2, 159, 2, 
/* out0016_had-eta8-phi22 */     3, 92, 4, 117, 4, 122, 2, 
/* out0017_had-eta8-phi23 */     2, 92, 4, 122, 4, 
/* out0018_had-eta9-phi22 */     5, 92, 2, 121, 2, 136, 2, 140, 6, 161, 4, 
/* out0019_had-eta9-phi23 */     5, 92, 2, 121, 6, 136, 4, 150, 2, 161, 4, 
/* out0020_had-eta9-phi24 */     1, 121, 2, 
/* out0021_had-eta10-phi22 */     7, 116, 2, 121, 2, 136, 2, 139, 2, 150, 4, 160, 2, 161, 4, 
/* out0022_had-eta10-phi23 */     4, 121, 4, 136, 4, 150, 4, 161, 4, 
/* out0023_had-eta6-phi22 */     6, 69, 2, 70, 2, 93, 2, 110, 6, 118, 6, 178, 3, 
/* out0024_had-eta6-phi23 */     3, 93, 6, 110, 6, 178, 3, 
/* out0025_had-eta6-phi24 */     1, 93, 2, 
/* out0026_had-eta7-phi22 */     4, 69, 4, 117, 2, 118, 4, 122, 2, 
/* out0027_had-eta7-phi23 */     3, 92, 2, 93, 4, 122, 6, 
/* out0028_had-eta7-phi24 */     1, 122, 2, 
/* out0029_had-eta4-phi22 */     4, 70, 2, 71, 6, 111, 2, 178, 1, 
/* out0030_had-eta4-phi23 */     4, 94, 4, 95, 4, 111, 4, 178, 1, 
/* out0031_had-eta5-phi22 */     5, 70, 6, 94, 2, 110, 2, 111, 4, 178, 4, 
/* out0032_had-eta5-phi23 */     5, 93, 2, 94, 8, 110, 2, 111, 6, 178, 4, 
/* out0033_had-eta5-phi24 */     1, 94, 2, 
/* out0034_had-eta3-phi22 */     3, 71, 6, 72, 6, 179, 1, 
/* out0035_had-eta3-phi23 */     2, 95, 10, 179, 1, 
/* out0036_had-eta3-phi24 */     1, 95, 2, 
/* out0037_had-eta1-phi23 */     2, 179, 2, 186, 5, 
/* out0038_had-eta2-phi23 */     3, 72, 2, 179, 1, 186, 3, 
/* out0039_had-eta2-phi24 */     0, 
/* out0040_had-eta15-phi16 */     6, 0, 2, 56, 2, 102, 2, 123, 2, 141, 2, 151, 2, 
/* out0041_had-eta15-phi17 */     6, 0, 2, 56, 2, 102, 2, 123, 2, 141, 2, 151, 2, 
/* out0042_had-eta15-phi18 */     6, 0, 2, 56, 2, 102, 2, 114, 2, 137, 2, 162, 2, 
/* out0043_had-eta15-phi19 */     6, 0, 2, 56, 2, 102, 2, 114, 2, 137, 2, 162, 2, 
/* out0044_had-eta16-phi16 */     5, 0, 2, 102, 2, 123, 2, 141, 2, 151, 2, 
/* out0045_had-eta16-phi17 */     6, 0, 2, 56, 2, 102, 2, 123, 2, 141, 2, 151, 2, 
/* out0046_had-eta16-phi18 */     3, 0, 2, 102, 2, 137, 2, 
/* out0047_had-eta16-phi19 */     3, 0, 2, 137, 2, 162, 2, 
/* out0048_had-eta11-phi19 */     2, 1, 2, 163, 2, 
/* out0049_had-eta12-phi18 */     1, 1, 2, 
/* out0050_had-eta12-phi19 */     3, 1, 2, 115, 2, 163, 2, 
/* out0051_had-eta12-phi20 */     4, 1, 2, 115, 2, 138, 4, 163, 4, 
/* out0052_had-eta13-phi18 */     1, 1, 2, 
/* out0053_had-eta13-phi19 */     5, 1, 2, 115, 2, 138, 2, 162, 2, 163, 2, 
/* out0054_had-eta13-phi20 */     4, 1, 2, 115, 2, 138, 2, 163, 2, 
/* out0055_had-eta14-phi19 */     5, 1, 2, 56, 2, 114, 2, 137, 2, 162, 2, 
/* out0056_had-eta9-phi19 */     1, 2, 2, 
/* out0057_had-eta9-phi20 */     3, 2, 4, 116, 2, 164, 2, 
/* out0058_had-eta9-phi21 */     4, 2, 2, 116, 4, 140, 8, 164, 2, 
/* out0059_had-eta10-phi19 */     1, 2, 2, 
/* out0060_had-eta10-phi20 */     4, 2, 2, 116, 2, 139, 2, 164, 4, 
/* out0061_had-eta10-phi21 */     4, 2, 2, 116, 4, 139, 4, 164, 4, 
/* out0062_had-eta11-phi20 */     5, 2, 2, 115, 2, 139, 2, 163, 2, 164, 2, 
/* out0063_had-eta7-phi20 */     0, 
/* out0064_had-eta7-phi21 */     3, 69, 6, 117, 4, 118, 2, 
/* out0065_had-eta8-phi20 */     0, 
/* out0066_had-eta8-phi21 */     2, 117, 6, 140, 2, 
/* out0067_had-eta5-phi21 */     2, 70, 4, 176, 4, 
/* out0068_had-eta6-phi21 */     3, 69, 4, 118, 4, 176, 2, 
/* out0069_had-eta3-phi21 */     3, 71, 2, 173, 1, 177, 1, 
/* out0070_had-eta4-phi21 */     4, 70, 2, 71, 2, 172, 8, 176, 2, 
/* out0071_had-eta2-phi21 */     3, 72, 2, 173, 1, 177, 1, 
/* out0072_had-eta2-phi22 */     3, 72, 6, 179, 1, 186, 3, 
/* out0073_had-eta1-phi22 */     2, 179, 2, 186, 5, 
/* out0074_had-eta16-phi1 */     2, 33, 2, 57, 2, 
/* out0075_had-eta16-phi2 */     2, 33, 2, 57, 2, 
/* out0076_had-eta16-phi3 */     0, 
/* out0077_had-eta16-phi4 */     0, 
/* out0078_had-eta17-phi1 */     1, 57, 2, 
/* out0079_had-eta17-phi2 */     0, 
/* out0080_had-eta17-phi3 */     0, 
/* out0081_had-eta17-phi4 */     0, 
/* out0082_had-eta16-phi7 */     0, 
/* out0083_had-eta16-phi8 */     0, 
/* out0084_had-eta16-phi9 */     0, 
/* out0085_had-eta16-phi10 */     1, 145, 2, 
/* out0086_had-eta17-phi6 */     0, 
/* out0087_had-eta17-phi8 */     0, 
/* out0088_had-eta17-phi9 */     0, 
/* out0089_had-eta17-phi10 */     0, 
/* out0090_had-eta14-phi12 */     2, 152, 2, 166, 2, 
/* out0091_had-eta14-phi13 */     2, 152, 2, 166, 2, 
/* out0092_had-eta14-phi14 */     3, 142, 2, 153, 2, 166, 2, 
/* out0093_had-eta15-phi12 */     2, 145, 2, 152, 2, 
/* out0094_had-eta15-phi13 */     2, 152, 2, 166, 2, 
/* out0095_had-eta15-phi14 */     3, 152, 2, 165, 2, 166, 2, 
/* out0096_had-eta16-phi12 */     1, 152, 2, 
/* out0097_had-eta16-phi13 */     2, 152, 2, 165, 2, 
/* out0098_had-eta12-phi15 */     5, 58, 2, 103, 2, 124, 4, 142, 4, 153, 2, 
/* out0099_had-eta12-phi16 */     3, 58, 2, 103, 2, 124, 2, 
/* out0100_had-eta12-phi17 */     2, 58, 2, 103, 2, 
/* out0101_had-eta13-phi15 */     4, 103, 2, 124, 2, 142, 2, 153, 2, 
/* out0102_had-eta13-phi16 */     5, 58, 2, 103, 2, 124, 2, 142, 2, 153, 2, 
/* out0103_had-eta13-phi17 */     2, 58, 2, 103, 2, 
/* out0104_had-eta14-phi15 */     3, 123, 2, 142, 2, 153, 2, 
/* out0105_had-eta14-phi16 */     4, 103, 2, 123, 2, 141, 2, 153, 2, 
/* out0106_had-eta9-phi17 */     0, 
/* out0107_had-eta9-phi18 */     0, 
/* out0108_had-eta10-phi16 */     2, 60, 2, 104, 2, 
/* out0109_had-eta10-phi17 */     0, 
/* out0110_had-eta10-phi18 */     0, 
/* out0111_had-eta11-phi17 */     1, 58, 2, 
/* out0112_had-eta11-phi18 */     0, 
/* out0113_had-eta7-phi18 */     2, 3, 2, 174, 2, 
/* out0114_had-eta7-phi19 */     1, 174, 2, 
/* out0115_had-eta8-phi18 */     1, 174, 2, 
/* out0116_had-eta8-phi19 */     1, 174, 2, 
/* out0117_had-eta5-phi19 */     4, 22, 4, 80, 4, 112, 8, 174, 2, 
/* out0118_had-eta5-phi20 */     1, 176, 4, 
/* out0119_had-eta6-phi19 */     2, 22, 2, 174, 2, 
/* out0120_had-eta6-phi20 */     1, 176, 2, 
/* out0121_had-eta4-phi19 */     4, 23, 8, 81, 6, 112, 4, 175, 1, 
/* out0122_had-eta4-phi20 */     3, 23, 2, 172, 8, 176, 2, 
/* out0123_had-eta2-phi20 */     4, 24, 6, 25, 4, 173, 1, 177, 1, 
/* out0124_had-eta3-phi20 */     3, 24, 4, 173, 1, 177, 1, 
/* out0125_had-eta1-phi20 */     4, 25, 10, 28, 2, 173, 2, 177, 1, 
/* out0126_had-eta1-phi21 */     2, 173, 2, 177, 1, 
/* out0127_had-eta0-phi21 */     2, 173, 2, 177, 2, 
/* out0128_had-eta0-phi22 */     2, 179, 2, 187, 8, 
/* out0129_had-eta12-phi1 */     2, 34, 2, 59, 2, 
/* out0130_had-eta12-phi2 */     1, 34, 2, 
/* out0131_had-eta13-phi1 */     2, 34, 2, 59, 2, 
/* out0132_had-eta13-phi2 */     0, 
/* out0133_had-eta13-phi3 */     0, 
/* out0134_had-eta14-phi1 */     1, 59, 2, 
/* out0135_had-eta14-phi2 */     0, 
/* out0136_had-eta14-phi3 */     0, 
/* out0137_had-eta13-phi4 */     0, 
/* out0138_had-eta13-phi5 */     0, 
/* out0139_had-eta13-phi6 */     0, 
/* out0140_had-eta13-phi7 */     0, 
/* out0141_had-eta14-phi4 */     0, 
/* out0142_had-eta14-phi5 */     0, 
/* out0143_had-eta14-phi6 */     0, 
/* out0144_had-eta14-phi7 */     0, 
/* out0145_had-eta12-phi9 */     0, 
/* out0146_had-eta12-phi10 */     1, 146, 2, 
/* out0147_had-eta13-phi8 */     0, 
/* out0148_had-eta13-phi9 */     0, 
/* out0149_had-eta13-phi10 */     1, 146, 2, 
/* out0150_had-eta14-phi8 */     0, 
/* out0151_had-eta14-phi9 */     0, 
/* out0152_had-eta14-phi10 */     1, 145, 2, 
/* out0153_had-eta11-phi12 */     3, 154, 2, 156, 2, 167, 2, 
/* out0154_had-eta11-phi13 */     4, 143, 2, 155, 2, 156, 2, 167, 4, 
/* out0155_had-eta12-phi11 */     2, 146, 4, 154, 2, 
/* out0156_had-eta12-phi12 */     3, 146, 2, 154, 4, 167, 2, 
/* out0157_had-eta12-phi13 */     2, 154, 2, 167, 4, 
/* out0158_had-eta12-phi14 */     4, 124, 2, 142, 2, 153, 2, 155, 2, 
/* out0159_had-eta13-phi12 */     2, 154, 2, 166, 2, 
/* out0160_had-eta13-phi13 */     2, 154, 2, 166, 2, 
/* out0161_had-eta9-phi14 */     6, 60, 2, 104, 2, 125, 2, 126, 2, 144, 8, 157, 6, 
/* out0162_had-eta9-phi15 */     2, 60, 4, 104, 2, 
/* out0163_had-eta9-phi16 */     2, 60, 2, 104, 2, 
/* out0164_had-eta10-phi14 */     6, 60, 2, 104, 2, 125, 4, 143, 4, 155, 4, 157, 2, 
/* out0165_had-eta10-phi15 */     5, 60, 2, 104, 4, 125, 4, 143, 2, 155, 2, 
/* out0166_had-eta11-phi14 */     4, 125, 2, 143, 4, 155, 4, 167, 2, 
/* out0167_had-eta11-phi15 */     6, 58, 2, 104, 2, 124, 2, 125, 2, 143, 2, 155, 2, 
/* out0168_had-eta7-phi16 */     0, 
/* out0169_had-eta7-phi17 */     1, 3, 2, 
/* out0170_had-eta8-phi15 */     1, 60, 2, 
/* out0171_had-eta8-phi16 */     0, 
/* out0172_had-eta8-phi17 */     0, 
/* out0173_had-eta5-phi17 */     3, 3, 2, 4, 4, 113, 4, 
/* out0174_had-eta5-phi18 */     6, 3, 2, 22, 6, 80, 8, 112, 2, 113, 4, 174, 2, 
/* out0175_had-eta6-phi17 */     1, 3, 4, 
/* out0176_had-eta6-phi18 */     4, 3, 4, 22, 2, 80, 2, 174, 2, 
/* out0177_had-eta4-phi18 */     8, 22, 2, 23, 2, 80, 2, 81, 2, 82, 4, 112, 2, 113, 4, 175, 1, 
/* out0178_had-eta2-phi19 */     6, 12, 2, 24, 4, 26, 2, 27, 6, 175, 1, 190, 6, 
/* out0179_had-eta3-phi18 */     5, 11, 4, 26, 6, 81, 2, 82, 2, 175, 1, 
/* out0180_had-eta3-phi19 */     5, 23, 4, 24, 2, 26, 2, 81, 6, 175, 1, 
/* out0181_had-eta1-phi19 */     8, 12, 2, 25, 2, 27, 6, 28, 8, 43, 2, 175, 2, 190, 2, 191, 1, 
/* out0182_had-eta0-phi20 */     3, 28, 2, 173, 2, 177, 2, 
/* out0183_had-eta9-phi1 */     2, 35, 2, 61, 2, 
/* out0184_had-eta9-phi2 */     0, 
/* out0185_had-eta10-phi0 */     2, 35, 2, 61, 4, 
/* out0186_had-eta10-phi1 */     2, 35, 2, 61, 2, 
/* out0187_had-eta10-phi2 */     0, 
/* out0188_had-eta11-phi0 */     3, 34, 2, 35, 2, 61, 2, 
/* out0189_had-eta11-phi1 */     2, 34, 2, 61, 2, 
/* out0190_had-eta11-phi2 */     0, 
/* out0191_had-eta10-phi3 */     0, 
/* out0192_had-eta10-phi4 */     2, 128, 2, 129, 2, 
/* out0193_had-eta10-phi5 */     3, 128, 2, 130, 2, 170, 4, 
/* out0194_had-eta11-phi3 */     1, 128, 2, 
/* out0195_had-eta11-phi4 */     1, 128, 4, 
/* out0196_had-eta11-phi5 */     1, 128, 4, 
/* out0197_had-eta12-phi4 */     1, 128, 2, 
/* out0198_had-eta12-phi5 */     0, 
/* out0199_had-eta10-phi6 */     2, 130, 2, 170, 6, 
/* out0200_had-eta10-phi7 */     1, 171, 6, 
/* out0201_had-eta10-phi8 */     1, 171, 4, 
/* out0202_had-eta11-phi6 */     2, 168, 4, 170, 2, 
/* out0203_had-eta11-phi7 */     1, 168, 4, 
/* out0204_had-eta11-phi8 */     0, 
/* out0205_had-eta12-phi7 */     1, 168, 4, 
/* out0206_had-eta12-phi8 */     0, 
/* out0207_had-eta9-phi9 */     0, 
/* out0208_had-eta9-phi10 */     0, 
/* out0209_had-eta10-phi9 */     0, 
/* out0210_had-eta10-phi10 */     1, 147, 4, 
/* out0211_had-eta10-phi11 */     2, 147, 4, 156, 2, 
/* out0212_had-eta11-phi9 */     0, 
/* out0213_had-eta11-phi10 */     1, 146, 2, 
/* out0214_had-eta11-phi11 */     2, 146, 2, 147, 2, 
/* out0215_had-eta8-phi12 */     0, 
/* out0216_had-eta8-phi13 */     1, 126, 4, 
/* out0217_had-eta9-phi11 */     1, 147, 4, 
/* out0218_had-eta9-phi12 */     2, 156, 2, 169, 4, 
/* out0219_had-eta9-phi13 */     4, 126, 2, 144, 6, 157, 6, 169, 4, 
/* out0220_had-eta10-phi12 */     3, 147, 2, 156, 4, 169, 4, 
/* out0221_had-eta7-phi13 */     1, 127, 10, 
/* out0222_had-eta7-phi14 */     2, 126, 2, 127, 6, 
/* out0223_had-eta7-phi15 */     0, 
/* out0224_had-eta8-phi14 */     2, 126, 6, 144, 2, 
/* out0225_had-eta5-phi15 */     0, 
/* out0226_had-eta5-phi16 */     1, 4, 2, 
/* out0227_had-eta6-phi15 */     0, 
/* out0228_had-eta6-phi16 */     0, 
/* out0229_had-eta4-phi16 */     3, 4, 4, 5, 2, 36, 2, 
/* out0230_had-eta4-phi17 */     3, 4, 6, 82, 6, 113, 4, 
/* out0231_had-eta3-phi17 */     5, 5, 2, 11, 4, 36, 2, 82, 4, 84, 10, 
/* out0232_had-eta1-phi18 */     9, 12, 8, 27, 2, 29, 4, 38, 8, 42, 2, 43, 12, 175, 2, 190, 2, 191, 1, 
/* out0233_had-eta2-phi18 */     8, 11, 4, 12, 4, 26, 6, 27, 2, 29, 4, 42, 6, 175, 1, 190, 6, 
/* out0234_had-eta0-phi19 */     3, 28, 4, 175, 2, 191, 4, 
/* out0235_had-eta7-phi0 */     2, 83, 2, 85, 2, 
/* out0236_had-eta7-phi1 */     1, 83, 2, 
/* out0237_had-eta7-phi2 */     1, 131, 2, 
/* out0238_had-eta8-phi0 */     1, 83, 4, 
/* out0239_had-eta8-phi1 */     1, 83, 4, 
/* out0240_had-eta8-phi2 */     0, 
/* out0241_had-eta7-phi3 */     1, 131, 8, 
/* out0242_had-eta8-phi3 */     2, 129, 2, 131, 4, 
/* out0243_had-eta8-phi4 */     3, 44, 4, 129, 4, 132, 2, 
/* out0244_had-eta9-phi3 */     1, 129, 4, 
/* out0245_had-eta9-phi4 */     1, 129, 4, 
/* out0246_had-eta8-phi5 */     3, 44, 4, 130, 2, 132, 4, 
/* out0247_had-eta8-phi6 */     2, 130, 2, 133, 4, 
/* out0248_had-eta9-phi5 */     2, 130, 4, 170, 2, 
/* out0249_had-eta9-phi6 */     2, 130, 4, 170, 2, 
/* out0250_had-eta7-phi8 */     0, 
/* out0251_had-eta8-phi7 */     1, 133, 2, 
/* out0252_had-eta8-phi8 */     0, 
/* out0253_had-eta8-phi9 */     0, 
/* out0254_had-eta9-phi7 */     1, 171, 4, 
/* out0255_had-eta9-phi8 */     1, 171, 2, 
/* out0256_had-eta7-phi9 */     0, 
/* out0257_had-eta7-phi10 */     0, 
/* out0258_had-eta7-phi11 */     0, 
/* out0259_had-eta8-phi10 */     0, 
/* out0260_had-eta8-phi11 */     0, 
/* out0261_had-eta6-phi11 */     1, 108, 6, 
/* out0262_had-eta6-phi12 */     0, 
/* out0263_had-eta6-phi13 */     0, 
/* out0264_had-eta7-phi12 */     0, 
/* out0265_had-eta5-phi13 */     0, 
/* out0266_had-eta5-phi14 */     0, 
/* out0267_had-eta6-phi14 */     0, 
/* out0268_had-eta4-phi14 */     0, 
/* out0269_had-eta4-phi15 */     0, 
/* out0270_had-eta2-phi16 */     6, 5, 2, 6, 6, 13, 2, 36, 2, 37, 2, 39, 8, 
/* out0271_had-eta3-phi15 */     1, 5, 2, 
/* out0272_had-eta3-phi16 */     3, 5, 8, 36, 10, 84, 2, 
/* out0273_had-eta1-phi17 */     8, 13, 8, 14, 2, 29, 4, 37, 2, 38, 8, 40, 6, 42, 2, 45, 12, 
/* out0274_had-eta2-phi17 */     6, 11, 4, 13, 4, 29, 4, 37, 12, 42, 6, 84, 4, 
/* out0275_had-eta5-phi0 */     2, 85, 2, 86, 6, 
/* out0276_had-eta5-phi1 */     0, 
/* out0277_had-eta6-phi0 */     1, 85, 8, 
/* out0278_had-eta6-phi1 */     1, 85, 2, 
/* out0279_had-eta5-phi2 */     0, 
/* out0280_had-eta6-phi2 */     0, 
/* out0281_had-eta6-phi3 */     1, 46, 4, 
/* out0282_had-eta6-phi4 */     2, 46, 6, 182, 3, 
/* out0283_had-eta6-phi5 */     2, 73, 6, 182, 3, 
/* out0284_had-eta7-phi4 */     3, 44, 4, 131, 2, 132, 4, 
/* out0285_had-eta7-phi5 */     3, 44, 4, 73, 2, 132, 6, 
/* out0286_had-eta6-phi6 */     3, 73, 6, 87, 6, 96, 2, 
/* out0287_had-eta6-phi7 */     1, 87, 4, 
/* out0288_had-eta7-phi6 */     2, 73, 2, 133, 6, 
/* out0289_had-eta7-phi7 */     1, 133, 4, 
/* out0290_had-eta5-phi8 */     2, 89, 2, 184, 3, 
/* out0291_had-eta5-phi9 */     1, 184, 3, 
/* out0292_had-eta6-phi8 */     1, 184, 1, 
/* out0293_had-eta6-phi9 */     1, 184, 1, 
/* out0294_had-eta5-phi10 */     2, 108, 2, 109, 2, 
/* out0295_had-eta5-phi11 */     2, 108, 2, 109, 4, 
/* out0296_had-eta6-phi10 */     1, 108, 6, 
/* out0297_had-eta4-phi12 */     0, 
/* out0298_had-eta4-phi13 */     0, 
/* out0299_had-eta5-phi12 */     0, 
/* out0300_had-eta3-phi13 */     0, 
/* out0301_had-eta3-phi14 */     0, 
/* out0302_had-eta2-phi14 */     0, 
/* out0303_had-eta2-phi15 */     2, 6, 6, 39, 6, 
/* out0304_had-eta1-phi15 */     3, 6, 2, 7, 10, 41, 10, 
/* out0305_had-eta1-phi16 */     8, 6, 2, 7, 2, 13, 2, 14, 6, 39, 2, 40, 10, 41, 4, 45, 2, 
/* out0306_had-eta0-phi16 */     2, 14, 6, 47, 10, 
/* out0307_had-eta3-phi0 */     1, 88, 10, 
/* out0308_had-eta3-phi1 */     0, 
/* out0309_had-eta4-phi0 */     2, 86, 6, 88, 4, 
/* out0310_had-eta4-phi1 */     0, 
/* out0311_had-eta4-phi2 */     0, 
/* out0312_had-eta4-phi3 */     1, 48, 8, 
/* out0313_had-eta4-phi4 */     6, 15, 2, 16, 4, 48, 2, 90, 2, 106, 2, 182, 1, 
/* out0314_had-eta5-phi3 */     2, 46, 2, 48, 4, 
/* out0315_had-eta5-phi4 */     4, 15, 4, 46, 4, 48, 2, 182, 4, 
/* out0316_had-eta4-phi5 */     11, 15, 4, 17, 2, 50, 2, 62, 6, 63, 2, 75, 4, 90, 4, 97, 6, 105, 2, 106, 6, 182, 1, 
/* out0317_had-eta4-phi6 */     14, 8, 6, 17, 2, 50, 2, 62, 6, 64, 2, 74, 4, 75, 4, 76, 2, 89, 2, 96, 2, 97, 6, 98, 2, 105, 2, 107, 6, 
/* out0318_had-eta5-phi5 */     4, 15, 6, 62, 2, 105, 6, 182, 4, 
/* out0319_had-eta5-phi6 */     5, 62, 2, 74, 6, 87, 4, 96, 8, 105, 6, 
/* out0320_had-eta4-phi7 */     7, 8, 2, 74, 2, 76, 6, 89, 6, 91, 2, 98, 8, 107, 2, 
/* out0321_had-eta4-phi8 */     4, 89, 2, 91, 2, 98, 2, 184, 4, 
/* out0322_had-eta5-phi7 */     4, 74, 4, 87, 2, 89, 4, 96, 4, 
/* out0323_had-eta4-phi9 */     1, 184, 4, 
/* out0324_had-eta4-phi10 */     1, 109, 4, 
/* out0325_had-eta3-phi10 */     0, 
/* out0326_had-eta3-phi11 */     0, 
/* out0327_had-eta4-phi11 */     1, 109, 6, 
/* out0328_had-eta3-phi12 */     0, 
/* out0329_had-eta2-phi13 */     0, 
/* out0330_had-eta1-phi14 */     0, 
/* out0331_had-eta0-phi15 */     2, 7, 4, 41, 2, 
/* out0332_had-eta2-phi0 */     0, 
/* out0333_had-eta2-phi1 */     0, 
/* out0334_had-eta2-phi2 */     1, 51, 8, 
/* out0335_had-eta3-phi2 */     1, 49, 4, 
/* out0336_had-eta3-phi3 */     2, 16, 2, 49, 10, 
/* out0337_had-eta3-phi4 */     7, 16, 8, 63, 4, 77, 2, 90, 2, 99, 4, 106, 2, 183, 1, 
/* out0338_had-eta3-phi5 */     14, 16, 2, 17, 6, 19, 2, 30, 6, 50, 6, 52, 2, 63, 10, 75, 4, 77, 8, 90, 8, 97, 2, 99, 12, 106, 6, 183, 1, 
/* out0339_had-eta3-phi6 */     11, 8, 6, 17, 6, 30, 8, 50, 6, 64, 10, 75, 4, 76, 2, 78, 6, 97, 2, 100, 12, 107, 6, 
/* out0340_had-eta3-phi7 */     11, 8, 2, 9, 4, 64, 4, 76, 6, 78, 2, 79, 4, 91, 6, 98, 4, 100, 2, 101, 8, 107, 2, 
/* out0341_had-eta3-phi8 */     4, 79, 2, 91, 6, 101, 6, 185, 1, 
/* out0342_had-eta2-phi9 */     2, 185, 1, 188, 6, 
/* out0343_had-eta3-phi9 */     1, 185, 1, 
/* out0344_had-eta2-phi10 */     1, 180, 4, 
/* out0345_had-eta2-phi11 */     1, 180, 4, 
/* out0346_had-eta1-phi12 */     0, 
/* out0347_had-eta2-phi12 */     0, 
/* out0348_had-eta1-phi13 */     0, 
/* out0349_had-eta0-phi13 */     0, 
/* out0350_had-eta0-phi14 */     0, 
/* out0351_had-eta1-phi0 */     0, 
/* out0352_had-eta1-phi1 */     0, 
/* out0353_had-eta1-phi2 */     2, 51, 2, 53, 10, 
/* out0354_had-eta2-phi3 */     3, 18, 8, 49, 2, 51, 4, 
/* out0355_had-eta2-phi4 */     8, 18, 6, 19, 4, 21, 2, 52, 2, 54, 2, 65, 10, 77, 2, 183, 1, 
/* out0356_had-eta2-phi5 */     5, 19, 10, 52, 12, 65, 4, 77, 4, 183, 1, 
/* out0357_had-eta2-phi6 */     6, 9, 2, 30, 2, 31, 12, 66, 4, 78, 6, 100, 2, 
/* out0358_had-eta2-phi7 */     7, 9, 10, 10, 2, 31, 2, 66, 10, 78, 2, 79, 6, 101, 2, 
/* out0359_had-eta2-phi8 */     3, 79, 4, 185, 1, 188, 6, 
/* out0360_had-eta1-phi9 */     3, 185, 1, 188, 2, 189, 1, 
/* out0361_had-eta1-phi10 */     1, 180, 4, 
/* out0362_had-eta1-phi11 */     1, 180, 4, 
/* out0363_had-eta0-phi1 */     0, 
/* out0364_had-eta0-phi2 */     1, 53, 4, 
/* out0365_had-eta1-phi3 */     5, 18, 2, 20, 12, 51, 2, 53, 2, 67, 2, 
/* out0366_had-eta1-phi4 */     7, 20, 2, 21, 10, 54, 10, 55, 2, 65, 2, 67, 12, 183, 2, 
/* out0367_had-eta1-phi5 */     3, 21, 4, 54, 4, 183, 2, 
/* out0368_had-eta1-phi6 */     2, 31, 2, 32, 4, 
/* out0369_had-eta1-phi7 */     4, 10, 8, 32, 10, 66, 2, 68, 12, 
/* out0370_had-eta1-phi8 */     5, 10, 6, 68, 2, 185, 1, 188, 2, 189, 1, 
/* out0371_had-eta0-phi9 */     2, 185, 2, 189, 4, 
/* out0372_had-eta0-phi10 */     1, 181, 7, 
/* out0373_had-eta16-phi20 */     2, 137, 2, 158, 2, 
/* out0374_had-eta16-phi21 */     2, 137, 2, 158, 2, 
/* out0375_had-eta17-phi19 */     0, 
/* out0376_had-eta17-phi20 */     1, 158, 2, 
/* out0377_had-eta17-phi21 */     1, 158, 2, 
/* out0378_had-eta17-phi22 */     1, 158, 2, 
/* out0379_had-eta12-phi21 */     3, 115, 2, 138, 2, 163, 2, 
/* out0380_had-eta13-phi21 */     3, 115, 2, 138, 2, 159, 2, 
/* out0381_had-eta14-phi20 */     3, 114, 2, 138, 2, 162, 2, 
/* out0382_had-eta11-phi21 */     5, 115, 2, 116, 2, 139, 4, 160, 2, 164, 2, 
/* out0383_had-eta16-phi14 */     3, 141, 2, 151, 2, 165, 2, 
/* out0384_had-eta16-phi15 */     4, 123, 2, 141, 2, 151, 2, 165, 2, 
/* out0385_had-eta17-phi13 */     1, 165, 2, 
/* out0386_had-eta17-phi14 */     1, 165, 2, 
/* out0387_had-eta17-phi15 */     1, 165, 2, 
/* out0388_had-eta17-phi16 */     1, 151, 2, 
/* out0389_had-eta17-phi17 */     0, 
/* out0390_had-eta14-phi17 */     2, 56, 2, 102, 2, 
/* out0391_had-eta14-phi18 */     3, 56, 2, 114, 2, 162, 2, 
/* out0392_had-eta14-phi0 */     1, 59, 2, 
/* out0393_had-eta15-phi0 */     2, 33, 2, 57, 2, 
/* out0394_had-eta15-phi1 */     2, 33, 2, 57, 2, 
/* out0395_had-eta15-phi2 */     2, 33, 2, 57, 2, 
/* out0396_had-eta16-phi0 */     2, 33, 2, 57, 2, 
/* out0397_had-eta15-phi4 */     0, 
/* out0398_had-eta15-phi5 */     0, 
/* out0399_had-eta15-phi6 */     0, 
/* out0400_had-eta16-phi5 */     0, 
/* out0401_had-eta16-phi6 */     0, 
/* out0402_had-eta14-phi11 */     1, 145, 2, 
/* out0403_had-eta15-phi9 */     1, 145, 2, 
/* out0404_had-eta15-phi10 */     1, 145, 2, 
/* out0405_had-eta15-phi11 */     2, 145, 2, 152, 2, 
/* out0406_had-eta16-phi11 */     1, 145, 2, 
/* out0407_had-eta13-phi14 */     4, 124, 2, 142, 2, 153, 2, 166, 2, 
/* out0408_had-eta11-phi16 */     2, 58, 2, 103, 2, 
/* out0409_had-eta12-phi-1 */     2, 34, 2, 59, 2, 
/* out0410_had-eta12-phi0 */     2, 34, 2, 59, 2, 
/* out0411_had-eta13-phi0 */     2, 34, 2, 59, 2, 
/* out0412_had-eta12-phi3 */     0, 
/* out0413_had-eta12-phi6 */     1, 168, 4, 
/* out0414_had-eta13-phi11 */     2, 146, 2, 154, 2, 
/* out0415_had-eta10-phi13 */     6, 125, 2, 143, 2, 156, 4, 157, 2, 167, 2, 169, 4, 
/* out0416_had-eta9-phi-1 */     1, 35, 2, 
/* out0417_had-eta9-phi0 */     3, 35, 4, 61, 2, 83, 2, 
/* out0418_had-eta0-phi18 */     3, 43, 2, 175, 2, 191, 4, 
/* out0419_had-eta7-phi-1 */     0, 
/* out0420_had-eta5-phi-1 */     1, 86, 2, 
/* out0421_had-eta0-phi17 */     3, 14, 2, 45, 2, 47, 6, 
/* out0422_had-eta3-phi-1 */     1, 88, 2, 
/* out0423_had-eta2-phi-1 */     0, 
/* out0424_had-eta0-phi0 */     0, 
/* out0425_had-eta1-phi-1 */     0, 
/* out0426_had-eta0-phi11 */     1, 181, 7, 
/* out0427_had-eta0-phi3 */     2, 20, 2, 55, 2, 
/* out0428_had-eta0-phi8 */     2, 185, 2, 189, 4, 
/* out0429_had-eta16-phi23 */     3, 134, 2, 148, 2, 158, 2, 
/* out0430_had-eta4-phi24 */     0, 
/* out0431_had-eta0-phi23 */     2, 179, 2, 187, 8, 
/* out0432_had-eta1-phi24 */     0, 
/* out0433_had-eta17-phi5 */     0, 
/* out0434_had-eta17-phi7 */     0, 
/* out0435_had-eta0-phi12 */     0, 
/* out0436_had-eta0-phi4 */     3, 55, 12, 67, 2, 183, 2, 
/* out0437_had-eta0-phi5 */     1, 183, 2, 
/* out0438_had-eta0-phi6 */     0, 
/* out0439_had-eta0-phi7 */     2, 32, 2, 68, 2, 
/* out0440_had-eta17-phi18 */     0, 
/* out0441_had-eta16-phi-1 */     1, 33, 2, 
/* out0442_had-eta17-phi11 */     0, 
/* out0443_had-eta4-phi-1 */     1, 86, 2, 
/* out0444_had-eta16-phi24 */     0, 
/* out0445_had-eta17-phi23 */     1, 158, 2, 
/* out0446_had-eta10-phi24 */     2, 136, 2, 150, 2, 
/* out0447_had-eta17-phi12 */     1, 165, 2, 
/* out0448_had-eta15-phi7 */     0, 
/* out0449_had-eta17-phi0 */     2, 33, 2, 57, 2, 
/* out0450_had-eta15-phi15 */     3, 123, 2, 141, 2, 151, 2, 
/* out0451_had-eta10-phi-1 */     2, 35, 2, 61, 2, 
/* out0452_had-eta8-phi-1 */     1, 83, 2, 
/* out0453_had-eta13-phi24 */     0, 
/* out0454_had-eta8-phi24 */     1, 92, 2, 
/* out0455_had-eta0-phi24 */     0, 
/* out0456_had-eta15-phi8 */     0, 
/* out0457_had-eta13-phi-1 */     1, 59, 2, 
/* out0458_had-eta15-phi3 */     0, 
/* out0459_had-eta6-phi-1 */     1, 85, 2, 
/* out0460_had-eta15-phi20 */     3, 114, 2, 137, 2, 162, 2, 
/* out0461_had-eta17-phi24 */     0, 
/* out0462_had-eta17-phi-1 */     0, 
/* out0463_had-eta11-phi-1 */     0, 
/* out0464_had-eta14-phi24 */     1, 119, 2, 
/* out0465_had-eta14-phi-1 */     0, 
/* out0466_had-eta15-phi-1 */     0, 
/* out0467_had-eta-2-phi0 */     0, 
/* out0468_had-eta-1-phi0 */     0, 
/* out0469_had-eta-2-phi1 */     0, 
/* out0470_had-eta-1-phi1 */     0, 
/* out0471_had-eta-2-phi2 */     0, 
/* out0472_had-eta-1-phi2 */     0, 
/* out0473_had-eta-2-phi3 */     0, 
/* out0474_had-eta-1-phi3 */     0, 
/* out0475_had-eta-2-phi4 */     0, 
/* out0476_had-eta-1-phi4 */     1, 183, 2, 
/* out0477_had-eta-2-phi5 */     0, 
/* out0478_had-eta-1-phi5 */     1, 183, 2, 
/* out0479_had-eta-2-phi6 */     0, 
/* out0480_had-eta-1-phi6 */     0, 
/* out0481_had-eta-2-phi7 */     0, 
/* out0482_had-eta-1-phi7 */     0, 
/* out0483_had-eta-2-phi8 */     1, 185, 1, 
/* out0484_had-eta-1-phi8 */     2, 185, 2, 189, 3, 
/* out0485_had-eta-2-phi9 */     1, 185, 1, 
/* out0486_had-eta-1-phi9 */     2, 185, 2, 189, 3, 
/* out0487_had-eta-2-phi10 */     0, 
/* out0488_had-eta-1-phi10 */     1, 181, 1, 
/* out0489_had-eta-2-phi11 */     0, 
/* out0490_had-eta-1-phi11 */     1, 181, 1, 
/* out0491_had-eta-2-phi12 */     0, 
/* out0492_had-eta-1-phi12 */     0, 
/* out0493_had-eta-2-phi13 */     0, 
/* out0494_had-eta-1-phi13 */     0, 
/* out0495_had-eta-2-phi14 */     0, 
/* out0496_had-eta-1-phi14 */     0, 
/* out0497_had-eta-2-phi15 */     0, 
/* out0498_had-eta-1-phi15 */     0, 
/* out0499_had-eta-2-phi16 */     0, 
/* out0500_had-eta-1-phi16 */     0, 
/* out0501_had-eta-2-phi17 */     0, 
/* out0502_had-eta-1-phi17 */     0, 
/* out0503_had-eta-2-phi18 */     0, 
/* out0504_had-eta-1-phi18 */     2, 175, 1, 191, 3, 
/* out0505_had-eta-2-phi19 */     0, 
/* out0506_had-eta-1-phi19 */     2, 175, 1, 191, 3, 
/* out0507_had-eta-2-phi20 */     1, 177, 1, 
/* out0508_had-eta-1-phi20 */     2, 173, 2, 177, 2, 
/* out0509_had-eta-2-phi21 */     1, 177, 1, 
/* out0510_had-eta-1-phi21 */     2, 173, 2, 177, 2, 
/* out0511_had-eta-2-phi22 */     0, 
/* out0512_had-eta-1-phi22 */     1, 179, 2, 
/* out0513_had-eta-2-phi23 */     0, 
/* out0514_had-eta-1-phi23 */     11792
};