parameter integer matrixH [0:1328] = {
/* num inputs = 80 (in0-in79) */
/* num outputs = 467 (out0-out466) */
/* max inputs per outputs = 6 */

/* out0_had-eta14-phi21 */     1, 71, 1, 
/* out1_had-eta14-phi22 */     2, 60, 1, 71, 1, 
/* out2_had-eta14-phi23 */     2, 60, 1, 71, 1, 
/* out3_had-eta15-phi21 */     2, 60, 1, 71, 1, 
/* out4_had-eta15-phi22 */     2, 60, 1, 71, 1, 
/* out5_had-eta15-phi23 */     1, 60, 1, 
/* out6_had-eta15-phi24 */     1, 60, 1, 
/* out7_had-eta16-phi22 */     2, 60, 1, 70, 1, 
/* out8_had-eta11-phi22 */     2, 62, 1, 72, 2, 
/* out9_had-eta11-phi23 */     3, 61, 1, 62, 1, 72, 1, 
/* out10_had-eta11-phi24 */     0, 
/* out11_had-eta12-phi22 */     2, 61, 2, 72, 2, 
/* out12_had-eta12-phi23 */     2, 61, 2, 72, 1, 
/* out13_had-eta12-phi24 */     1, 61, 1, 
/* out14_had-eta13-phi22 */     2, 61, 1, 71, 1, 
/* out15_had-eta13-phi23 */     2, 61, 1, 71, 1, 
/* out16_had-eta8-phi22 */     1, 34, 2, 
/* out17_had-eta8-phi23 */     1, 34, 2, 
/* out18_had-eta9-phi22 */     2, 34, 1, 73, 2, 
/* out19_had-eta9-phi23 */     3, 34, 1, 62, 1, 73, 2, 
/* out20_had-eta9-phi24 */     0, 
/* out21_had-eta10-phi22 */     3, 62, 2, 72, 1, 73, 2, 
/* out22_had-eta10-phi23 */     2, 62, 2, 73, 2, 
/* out23_had-eta6-phi22 */     1, 35, 1, 
/* out24_had-eta6-phi23 */     1, 35, 3, 
/* out25_had-eta6-phi24 */     1, 35, 1, 
/* out26_had-eta7-phi22 */     0, 
/* out27_had-eta7-phi23 */     2, 34, 1, 35, 2, 
/* out28_had-eta7-phi24 */     0, 
/* out29_had-eta4-phi22 */     0, 
/* out30_had-eta4-phi23 */     2, 36, 2, 37, 2, 
/* out31_had-eta5-phi22 */     1, 36, 1, 
/* out32_had-eta5-phi23 */     2, 35, 1, 36, 4, 
/* out33_had-eta5-phi24 */     1, 36, 1, 
/* out34_had-eta3-phi22 */     0, 
/* out35_had-eta3-phi23 */     1, 37, 5, 
/* out36_had-eta3-phi24 */     1, 37, 1, 
/* out37_had-eta1-phi23 */     0, 
/* out38_had-eta2-phi23 */     0, 
/* out39_had-eta2-phi24 */     0, 
/* out40_had-eta15-phi16 */     1, 63, 1, 
/* out41_had-eta15-phi17 */     1, 63, 1, 
/* out42_had-eta15-phi18 */     0, 
/* out43_had-eta15-phi19 */     0, 
/* out44_had-eta16-phi16 */     1, 63, 1, 
/* out45_had-eta16-phi17 */     1, 63, 1, 
/* out46_had-eta16-phi18 */     0, 
/* out47_had-eta16-phi19 */     0, 
/* out48_had-eta11-phi19 */     0, 
/* out49_had-eta12-phi18 */     0, 
/* out50_had-eta12-phi19 */     0, 
/* out51_had-eta12-phi20 */     0, 
/* out52_had-eta13-phi18 */     0, 
/* out53_had-eta13-phi19 */     0, 
/* out54_had-eta13-phi20 */     0, 
/* out55_had-eta14-phi19 */     0, 
/* out56_had-eta9-phi19 */     0, 
/* out57_had-eta9-phi20 */     0, 
/* out58_had-eta9-phi21 */     0, 
/* out59_had-eta10-phi19 */     0, 
/* out60_had-eta10-phi20 */     0, 
/* out61_had-eta10-phi21 */     0, 
/* out62_had-eta11-phi20 */     0, 
/* out63_had-eta7-phi20 */     1, 29, 2, 
/* out64_had-eta7-phi21 */     0, 
/* out65_had-eta8-phi20 */     1, 29, 1, 
/* out66_had-eta8-phi21 */     0, 
/* out67_had-eta5-phi21 */     2, 30, 1, 31, 1, 
/* out68_had-eta6-phi21 */     1, 30, 1, 
/* out69_had-eta3-phi21 */     1, 32, 4, 
/* out70_had-eta4-phi21 */     1, 31, 3, 
/* out71_had-eta2-phi21 */     1, 32, 2, 
/* out72_had-eta2-phi22 */     0, 
/* out73_had-eta1-phi22 */     0, 
/* out74_had-eta16-phi1 */     0, 
/* out75_had-eta16-phi2 */     0, 
/* out76_had-eta16-phi3 */     0, 
/* out77_had-eta16-phi4 */     1, 5, 1, 
/* out78_had-eta17-phi1 */     0, 
/* out79_had-eta17-phi2 */     0, 
/* out80_had-eta17-phi3 */     0, 
/* out81_had-eta17-phi4 */     0, 
/* out82_had-eta16-phi7 */     1, 5, 1, 
/* out83_had-eta16-phi8 */     1, 47, 1, 
/* out84_had-eta16-phi9 */     1, 47, 1, 
/* out85_had-eta16-phi10 */     4, 6, 1, 47, 1, 51, 1, 74, 1, 
/* out86_had-eta17-phi6 */     1, 5, 1, 
/* out87_had-eta17-phi8 */     0, 
/* out88_had-eta17-phi9 */     0, 
/* out89_had-eta17-phi10 */     0, 
/* out90_had-eta14-phi12 */     2, 11, 1, 64, 1, 
/* out91_had-eta14-phi13 */     2, 11, 1, 64, 1, 
/* out92_had-eta14-phi14 */     1, 65, 1, 
/* out93_had-eta15-phi12 */     5, 11, 1, 18, 1, 51, 1, 64, 1, 74, 1, 
/* out94_had-eta15-phi13 */     3, 11, 1, 18, 1, 64, 1, 
/* out95_had-eta15-phi14 */     3, 11, 1, 18, 1, 64, 1, 
/* out96_had-eta16-phi12 */     4, 6, 1, 11, 1, 18, 1, 64, 1, 
/* out97_had-eta16-phi13 */     3, 11, 1, 18, 1, 64, 1, 
/* out98_had-eta12-phi15 */     1, 65, 1, 
/* out99_had-eta12-phi16 */     0, 
/* out100_had-eta12-phi17 */     0, 
/* out101_had-eta13-phi15 */     1, 65, 1, 
/* out102_had-eta13-phi16 */     1, 65, 1, 
/* out103_had-eta13-phi17 */     0, 
/* out104_had-eta14-phi15 */     1, 65, 1, 
/* out105_had-eta14-phi16 */     1, 65, 1, 
/* out106_had-eta9-phi17 */     0, 
/* out107_had-eta9-phi18 */     0, 
/* out108_had-eta10-phi16 */     0, 
/* out109_had-eta10-phi17 */     0, 
/* out110_had-eta10-phi18 */     0, 
/* out111_had-eta11-phi17 */     0, 
/* out112_had-eta11-phi18 */     0, 
/* out113_had-eta7-phi18 */     1, 0, 1, 
/* out114_had-eta7-phi19 */     1, 29, 3, 
/* out115_had-eta8-phi18 */     0, 
/* out116_had-eta8-phi19 */     1, 29, 1, 
/* out117_had-eta5-phi19 */     2, 30, 1, 38, 4, 
/* out118_had-eta5-phi20 */     1, 30, 3, 
/* out119_had-eta6-phi19 */     1, 29, 1, 
/* out120_had-eta6-phi20 */     1, 30, 2, 
/* out121_had-eta4-phi19 */     2, 14, 2, 38, 2, 
/* out122_had-eta4-phi20 */     1, 31, 3, 
/* out123_had-eta2-phi20 */     2, 16, 2, 32, 1, 
/* out124_had-eta3-phi20 */     3, 15, 1, 31, 1, 32, 1, 
/* out125_had-eta1-phi20 */     2, 16, 1, 17, 4, 
/* out126_had-eta1-phi21 */     0, 
/* out127_had-eta0-phi21 */     0, 
/* out128_had-eta0-phi22 */     0, 
/* out129_had-eta12-phi1 */     0, 
/* out130_had-eta12-phi2 */     0, 
/* out131_had-eta13-phi1 */     0, 
/* out132_had-eta13-phi2 */     0, 
/* out133_had-eta13-phi3 */     1, 7, 1, 
/* out134_had-eta14-phi1 */     0, 
/* out135_had-eta14-phi2 */     0, 
/* out136_had-eta14-phi3 */     1, 7, 1, 
/* out137_had-eta13-phi4 */     2, 7, 1, 52, 1, 
/* out138_had-eta13-phi5 */     2, 7, 1, 52, 1, 
/* out139_had-eta13-phi6 */     1, 52, 2, 
/* out140_had-eta13-phi7 */     0, 
/* out141_had-eta14-phi4 */     2, 7, 1, 52, 1, 
/* out142_had-eta14-phi5 */     1, 52, 1, 
/* out143_had-eta14-phi6 */     1, 52, 1, 
/* out144_had-eta14-phi7 */     0, 
/* out145_had-eta12-phi9 */     2, 8, 1, 48, 1, 
/* out146_had-eta12-phi10 */     5, 8, 1, 48, 1, 49, 1, 53, 1, 75, 1, 
/* out147_had-eta13-phi8 */     0, 
/* out148_had-eta13-phi9 */     1, 48, 1, 
/* out149_had-eta13-phi10 */     4, 8, 1, 48, 1, 53, 1, 75, 1, 
/* out150_had-eta14-phi8 */     0, 
/* out151_had-eta14-phi9 */     1, 48, 1, 
/* out152_had-eta14-phi10 */     4, 6, 1, 48, 1, 51, 1, 74, 1, 
/* out153_had-eta11-phi12 */     4, 12, 1, 19, 1, 66, 1, 68, 1, 
/* out154_had-eta11-phi13 */     4, 12, 1, 19, 1, 67, 1, 68, 1, 
/* out155_had-eta12-phi11 */     6, 8, 1, 12, 1, 19, 1, 53, 2, 66, 1, 75, 2, 
/* out156_had-eta12-phi12 */     6, 8, 1, 12, 1, 19, 1, 53, 1, 66, 2, 75, 1, 
/* out157_had-eta12-phi13 */     3, 12, 1, 19, 1, 66, 1, 
/* out158_had-eta12-phi14 */     4, 12, 1, 19, 1, 65, 1, 67, 1, 
/* out159_had-eta13-phi12 */     4, 12, 1, 19, 1, 66, 1, 75, 1, 
/* out160_had-eta13-phi13 */     3, 12, 1, 19, 1, 66, 1, 
/* out161_had-eta9-phi14 */     1, 69, 3, 
/* out162_had-eta9-phi15 */     0, 
/* out163_had-eta9-phi16 */     0, 
/* out164_had-eta10-phi14 */     2, 67, 2, 69, 1, 
/* out165_had-eta10-phi15 */     1, 67, 1, 
/* out166_had-eta11-phi14 */     1, 67, 2, 
/* out167_had-eta11-phi15 */     1, 67, 1, 
/* out168_had-eta7-phi16 */     0, 
/* out169_had-eta7-phi17 */     1, 0, 1, 
/* out170_had-eta8-phi15 */     0, 
/* out171_had-eta8-phi16 */     0, 
/* out172_had-eta8-phi17 */     0, 
/* out173_had-eta5-phi17 */     5, 0, 1, 1, 2, 21, 2, 25, 1, 39, 2, 
/* out174_had-eta5-phi18 */     5, 0, 1, 14, 1, 25, 1, 38, 1, 39, 2, 
/* out175_had-eta6-phi17 */     1, 0, 2, 
/* out176_had-eta6-phi18 */     1, 0, 2, 
/* out177_had-eta4-phi18 */     5, 14, 4, 22, 1, 25, 3, 38, 1, 39, 2, 
/* out178_had-eta2-phi19 */     3, 15, 2, 16, 3, 23, 1, 
/* out179_had-eta3-phi18 */     3, 14, 1, 15, 1, 22, 3, 
/* out180_had-eta3-phi19 */     1, 15, 4, 
/* out181_had-eta1-phi19 */     3, 16, 2, 17, 1, 24, 5, 
/* out182_had-eta0-phi20 */     1, 17, 2, 
/* out183_had-eta9-phi1 */     0, 
/* out184_had-eta9-phi2 */     1, 9, 1, 
/* out185_had-eta10-phi0 */     0, 
/* out186_had-eta10-phi1 */     0, 
/* out187_had-eta10-phi2 */     1, 9, 1, 
/* out188_had-eta11-phi0 */     0, 
/* out189_had-eta11-phi1 */     0, 
/* out190_had-eta11-phi2 */     1, 9, 1, 
/* out191_had-eta10-phi3 */     2, 9, 1, 57, 1, 
/* out192_had-eta10-phi4 */     4, 9, 1, 41, 2, 54, 1, 57, 2, 
/* out193_had-eta10-phi5 */     3, 41, 2, 58, 2, 78, 2, 
/* out194_had-eta11-phi3 */     2, 9, 1, 54, 1, 
/* out195_had-eta11-phi4 */     1, 54, 2, 
/* out196_had-eta11-phi5 */     2, 40, 2, 54, 2, 
/* out197_had-eta12-phi4 */     2, 7, 1, 54, 1, 
/* out198_had-eta12-phi5 */     3, 7, 1, 40, 1, 54, 1, 
/* out199_had-eta10-phi6 */     5, 40, 1, 42, 2, 55, 1, 58, 2, 78, 3, 
/* out200_had-eta10-phi7 */     4, 42, 2, 55, 1, 59, 2, 79, 3, 
/* out201_had-eta10-phi8 */     2, 59, 1, 79, 2, 
/* out202_had-eta11-phi6 */     4, 40, 2, 55, 2, 76, 2, 78, 1, 
/* out203_had-eta11-phi7 */     2, 55, 2, 76, 2, 
/* out204_had-eta11-phi8 */     0, 
/* out205_had-eta12-phi7 */     2, 55, 1, 76, 2, 
/* out206_had-eta12-phi8 */     0, 
/* out207_had-eta9-phi9 */     0, 
/* out208_had-eta9-phi10 */     2, 10, 1, 50, 4, 
/* out209_had-eta10-phi9 */     0, 
/* out210_had-eta10-phi10 */     4, 10, 1, 49, 2, 56, 2, 77, 1, 
/* out211_had-eta10-phi11 */     6, 10, 1, 20, 1, 49, 1, 56, 2, 68, 1, 77, 2, 
/* out212_had-eta11-phi9 */     1, 49, 1, 
/* out213_had-eta11-phi10 */     4, 8, 1, 49, 2, 53, 1, 77, 1, 
/* out214_had-eta11-phi11 */     5, 8, 1, 49, 1, 53, 1, 56, 1, 77, 2, 
/* out215_had-eta8-phi12 */     1, 13, 1, 
/* out216_had-eta8-phi13 */     1, 13, 1, 
/* out217_had-eta9-phi11 */     6, 10, 2, 13, 1, 20, 1, 50, 3, 56, 2, 77, 1, 
/* out218_had-eta9-phi12 */     4, 10, 1, 13, 2, 20, 2, 68, 1, 
/* out219_had-eta9-phi13 */     3, 13, 1, 20, 1, 69, 3, 
/* out220_had-eta10-phi12 */     5, 13, 1, 20, 2, 56, 1, 68, 2, 77, 1, 
/* out221_had-eta7-phi13 */     0, 
/* out222_had-eta7-phi14 */     0, 
/* out223_had-eta7-phi15 */     0, 
/* out224_had-eta8-phi14 */     0, 
/* out225_had-eta5-phi15 */     0, 
/* out226_had-eta5-phi16 */     2, 1, 1, 21, 1, 
/* out227_had-eta6-phi15 */     0, 
/* out228_had-eta6-phi16 */     0, 
/* out229_had-eta4-phi16 */     3, 1, 2, 2, 1, 21, 2, 
/* out230_had-eta4-phi17 */     5, 1, 3, 21, 3, 22, 1, 25, 3, 39, 2, 
/* out231_had-eta3-phi17 */     3, 2, 1, 22, 3, 26, 5, 
/* out232_had-eta1-phi18 */     2, 23, 1, 24, 3, 
/* out233_had-eta2-phi18 */     1, 23, 6, 
/* out234_had-eta0-phi19 */     1, 17, 1, 
/* out235_had-eta7-phi0 */     0, 
/* out236_had-eta7-phi1 */     0, 
/* out237_had-eta7-phi2 */     0, 
/* out238_had-eta8-phi0 */     0, 
/* out239_had-eta8-phi1 */     0, 
/* out240_had-eta8-phi2 */     0, 
/* out241_had-eta7-phi3 */     1, 43, 1, 
/* out242_had-eta8-phi3 */     1, 43, 2, 
/* out243_had-eta8-phi4 */     1, 43, 3, 
/* out244_had-eta9-phi3 */     2, 9, 2, 57, 2, 
/* out245_had-eta9-phi4 */     2, 41, 2, 57, 3, 
/* out246_had-eta8-phi5 */     1, 44, 2, 
/* out247_had-eta8-phi6 */     1, 44, 3, 
/* out248_had-eta9-phi5 */     3, 41, 2, 58, 2, 78, 1, 
/* out249_had-eta9-phi6 */     3, 42, 2, 58, 2, 78, 1, 
/* out250_had-eta7-phi8 */     1, 45, 1, 
/* out251_had-eta8-phi7 */     1, 45, 3, 
/* out252_had-eta8-phi8 */     1, 45, 2, 
/* out253_had-eta8-phi9 */     0, 
/* out254_had-eta9-phi7 */     3, 42, 2, 59, 3, 79, 2, 
/* out255_had-eta9-phi8 */     2, 59, 2, 79, 1, 
/* out256_had-eta7-phi9 */     0, 
/* out257_had-eta7-phi10 */     1, 46, 4, 
/* out258_had-eta7-phi11 */     1, 46, 4, 
/* out259_had-eta8-phi10 */     2, 10, 1, 50, 1, 
/* out260_had-eta8-phi11 */     1, 10, 1, 
/* out261_had-eta6-phi11 */     0, 
/* out262_had-eta6-phi12 */     0, 
/* out263_had-eta6-phi13 */     0, 
/* out264_had-eta7-phi12 */     0, 
/* out265_had-eta5-phi13 */     0, 
/* out266_had-eta5-phi14 */     0, 
/* out267_had-eta6-phi14 */     0, 
/* out268_had-eta4-phi14 */     0, 
/* out269_had-eta4-phi15 */     0, 
/* out270_had-eta2-phi16 */     3, 2, 1, 3, 3, 27, 4, 
/* out271_had-eta3-phi15 */     1, 2, 1, 
/* out272_had-eta3-phi16 */     2, 2, 4, 26, 2, 
/* out273_had-eta1-phi17 */     0, 
/* out274_had-eta2-phi17 */     2, 26, 1, 27, 2, 
/* out275_had-eta5-phi0 */     0, 
/* out276_had-eta5-phi1 */     0, 
/* out277_had-eta6-phi0 */     0, 
/* out278_had-eta6-phi1 */     0, 
/* out279_had-eta5-phi2 */     0, 
/* out280_had-eta6-phi2 */     0, 
/* out281_had-eta6-phi3 */     0, 
/* out282_had-eta6-phi4 */     0, 
/* out283_had-eta6-phi5 */     0, 
/* out284_had-eta7-phi4 */     1, 43, 2, 
/* out285_had-eta7-phi5 */     1, 44, 1, 
/* out286_had-eta6-phi6 */     0, 
/* out287_had-eta6-phi7 */     0, 
/* out288_had-eta7-phi6 */     1, 44, 2, 
/* out289_had-eta7-phi7 */     1, 45, 2, 
/* out290_had-eta5-phi8 */     0, 
/* out291_had-eta5-phi9 */     0, 
/* out292_had-eta6-phi8 */     0, 
/* out293_had-eta6-phi9 */     0, 
/* out294_had-eta5-phi10 */     0, 
/* out295_had-eta5-phi11 */     0, 
/* out296_had-eta6-phi10 */     0, 
/* out297_had-eta4-phi12 */     0, 
/* out298_had-eta4-phi13 */     0, 
/* out299_had-eta5-phi12 */     0, 
/* out300_had-eta3-phi13 */     0, 
/* out301_had-eta3-phi14 */     0, 
/* out302_had-eta2-phi14 */     0, 
/* out303_had-eta2-phi15 */     1, 3, 3, 
/* out304_had-eta1-phi15 */     3, 3, 1, 4, 5, 28, 1, 
/* out305_had-eta1-phi16 */     4, 3, 1, 4, 1, 27, 2, 28, 5, 
/* out306_had-eta0-phi16 */     1, 28, 2, 
/* out307_had-eta3-phi0 */     0, 
/* out308_had-eta3-phi1 */     0, 
/* out309_had-eta4-phi0 */     0, 
/* out310_had-eta4-phi1 */     0, 
/* out311_had-eta4-phi2 */     0, 
/* out312_had-eta4-phi3 */     0, 
/* out313_had-eta4-phi4 */     1, 33, 1, 
/* out314_had-eta5-phi3 */     0, 
/* out315_had-eta5-phi4 */     0, 
/* out316_had-eta4-phi5 */     1, 33, 2, 
/* out317_had-eta4-phi6 */     0, 
/* out318_had-eta5-phi5 */     0, 
/* out319_had-eta5-phi6 */     0, 
/* out320_had-eta4-phi7 */     0, 
/* out321_had-eta4-phi8 */     0, 
/* out322_had-eta5-phi7 */     0, 
/* out323_had-eta4-phi9 */     0, 
/* out324_had-eta4-phi10 */     0, 
/* out325_had-eta3-phi10 */     0, 
/* out326_had-eta3-phi11 */     0, 
/* out327_had-eta4-phi11 */     0, 
/* out328_had-eta3-phi12 */     0, 
/* out329_had-eta2-phi13 */     0, 
/* out330_had-eta1-phi14 */     0, 
/* out331_had-eta0-phi15 */     1, 4, 2, 
/* out332_had-eta2-phi0 */     0, 
/* out333_had-eta2-phi1 */     0, 
/* out334_had-eta2-phi2 */     0, 
/* out335_had-eta3-phi2 */     0, 
/* out336_had-eta3-phi3 */     0, 
/* out337_had-eta3-phi4 */     1, 33, 1, 
/* out338_had-eta3-phi5 */     1, 33, 4, 
/* out339_had-eta3-phi6 */     0, 
/* out340_had-eta3-phi7 */     0, 
/* out341_had-eta3-phi8 */     0, 
/* out342_had-eta2-phi9 */     0, 
/* out343_had-eta3-phi9 */     0, 
/* out344_had-eta2-phi10 */     0, 
/* out345_had-eta2-phi11 */     0, 
/* out346_had-eta1-phi12 */     0, 
/* out347_had-eta2-phi12 */     0, 
/* out348_had-eta1-phi13 */     0, 
/* out349_had-eta0-phi13 */     0, 
/* out350_had-eta0-phi14 */     0, 
/* out351_had-eta1-phi0 */     0, 
/* out352_had-eta1-phi1 */     0, 
/* out353_had-eta1-phi2 */     0, 
/* out354_had-eta2-phi3 */     0, 
/* out355_had-eta2-phi4 */     0, 
/* out356_had-eta2-phi5 */     0, 
/* out357_had-eta2-phi6 */     0, 
/* out358_had-eta2-phi7 */     0, 
/* out359_had-eta2-phi8 */     0, 
/* out360_had-eta1-phi9 */     0, 
/* out361_had-eta1-phi10 */     0, 
/* out362_had-eta1-phi11 */     0, 
/* out363_had-eta0-phi1 */     0, 
/* out364_had-eta0-phi2 */     0, 
/* out365_had-eta1-phi3 */     0, 
/* out366_had-eta1-phi4 */     0, 
/* out367_had-eta1-phi5 */     0, 
/* out368_had-eta1-phi6 */     0, 
/* out369_had-eta1-phi7 */     0, 
/* out370_had-eta1-phi8 */     0, 
/* out371_had-eta0-phi9 */     0, 
/* out372_had-eta0-phi10 */     0, 
/* out373_had-eta16-phi20 */     1, 70, 1, 
/* out374_had-eta16-phi21 */     1, 70, 1, 
/* out375_had-eta17-phi19 */     0, 
/* out376_had-eta17-phi20 */     1, 70, 1, 
/* out377_had-eta17-phi21 */     1, 70, 1, 
/* out378_had-eta17-phi22 */     1, 70, 1, 
/* out379_had-eta12-phi21 */     0, 
/* out380_had-eta13-phi21 */     1, 71, 1, 
/* out381_had-eta14-phi20 */     0, 
/* out382_had-eta11-phi21 */     1, 72, 1, 
/* out383_had-eta16-phi14 */     3, 11, 1, 18, 1, 63, 1, 
/* out384_had-eta16-phi15 */     1, 63, 1, 
/* out385_had-eta17-phi13 */     0, 
/* out386_had-eta17-phi14 */     0, 
/* out387_had-eta17-phi15 */     0, 
/* out388_had-eta17-phi16 */     1, 63, 1, 
/* out389_had-eta17-phi17 */     0, 
/* out390_had-eta14-phi17 */     0, 
/* out391_had-eta14-phi18 */     0, 
/* out392_had-eta14-phi0 */     0, 
/* out393_had-eta15-phi0 */     0, 
/* out394_had-eta15-phi1 */     0, 
/* out395_had-eta15-phi2 */     0, 
/* out396_had-eta16-phi0 */     0, 
/* out397_had-eta15-phi4 */     1, 5, 1, 
/* out398_had-eta15-phi5 */     1, 5, 1, 
/* out399_had-eta15-phi6 */     1, 5, 1, 
/* out400_had-eta16-phi5 */     1, 5, 1, 
/* out401_had-eta16-phi6 */     1, 5, 1, 
/* out402_had-eta14-phi11 */     4, 6, 1, 48, 1, 51, 1, 74, 1, 
/* out403_had-eta15-phi9 */     4, 6, 1, 47, 2, 51, 1, 74, 1, 
/* out404_had-eta15-phi10 */     4, 6, 1, 47, 1, 51, 1, 74, 1, 
/* out405_had-eta15-phi11 */     4, 6, 1, 51, 1, 64, 1, 74, 1, 
/* out406_had-eta16-phi11 */     5, 6, 1, 18, 1, 47, 1, 51, 1, 74, 1, 
/* out407_had-eta13-phi14 */     1, 65, 1, 
/* out408_had-eta11-phi16 */     0, 
/* out409_had-eta12-phi-1 */     0, 
/* out410_had-eta12-phi0 */     0, 
/* out411_had-eta13-phi0 */     0, 
/* out412_had-eta12-phi3 */     1, 7, 1, 
/* out413_had-eta12-phi6 */     4, 40, 2, 52, 1, 55, 1, 76, 2, 
/* out414_had-eta13-phi11 */     5, 8, 1, 48, 1, 53, 1, 66, 1, 75, 2, 
/* out415_had-eta10-phi13 */     4, 13, 1, 20, 1, 68, 2, 69, 1, 
/* out416_had-eta9-phi-1 */     0, 
/* out417_had-eta9-phi0 */     0, 
/* out418_had-eta0-phi18 */     0, 
/* out419_had-eta7-phi-1 */     0, 
/* out420_had-eta5-phi-1 */     0, 
/* out421_had-eta0-phi17 */     0, 
/* out422_had-eta3-phi-1 */     0, 
/* out423_had-eta2-phi-1 */     0, 
/* out424_had-eta0-phi0 */     0, 
/* out425_had-eta1-phi-1 */     0, 
/* out426_had-eta0-phi11 */     0, 
/* out427_had-eta0-phi3 */     0, 
/* out428_had-eta0-phi8 */     0, 
/* out429_had-eta16-phi23 */     2, 60, 1, 70, 1, 
/* out430_had-eta4-phi24 */     0, 
/* out431_had-eta0-phi23 */     0, 
/* out432_had-eta1-phi24 */     0, 
/* out433_had-eta17-phi5 */     0, 
/* out434_had-eta17-phi7 */     0, 
/* out435_had-eta0-phi12 */     0, 
/* out436_had-eta0-phi4 */     0, 
/* out437_had-eta0-phi5 */     0, 
/* out438_had-eta0-phi6 */     0, 
/* out439_had-eta0-phi7 */     0, 
/* out440_had-eta17-phi18 */     0, 
/* out441_had-eta16-phi-1 */     0, 
/* out442_had-eta17-phi11 */     0, 
/* out443_had-eta4-phi-1 */     0, 
/* out444_had-eta16-phi24 */     0, 
/* out445_had-eta17-phi23 */     1, 70, 1, 
/* out446_had-eta10-phi24 */     1, 62, 1, 
/* out447_had-eta17-phi12 */     1, 18, 1, 
/* out448_had-eta15-phi7 */     0, 
/* out449_had-eta17-phi0 */     0, 
/* out450_had-eta15-phi15 */     1, 63, 1, 
/* out451_had-eta10-phi-1 */     0, 
/* out452_had-eta8-phi-1 */     0, 
/* out453_had-eta13-phi24 */     0, 
/* out454_had-eta8-phi24 */     1, 34, 1, 
/* out455_had-eta0-phi24 */     0, 
/* out456_had-eta15-phi8 */     1, 47, 1, 
/* out457_had-eta13-phi-1 */     0, 
/* out458_had-eta15-phi3 */     0, 
/* out459_had-eta6-phi-1 */     0, 
/* out460_had-eta15-phi20 */     0, 
/* out461_had-eta17-phi24 */     0, 
/* out462_had-eta17-phi-1 */     0, 
/* out463_had-eta11-phi-1 */     0, 
/* out464_had-eta14-phi24 */     0, 
/* out465_had-eta14-phi-1 */     0, 
/* out466_had-eta15-phi-1 */     0

};
