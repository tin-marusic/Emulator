parameter integer matrixH [0:2398] = {
/* num inputs = 161 (in0-in160) */
/* num outputs = 515(out0-out514) */
//* max inputs per outputs = 8 */
//* total number of input in adders 942 */

/* out0000_had-eta14-phi21 */     0, 
/* out0001_had-eta14-phi22 */     1, 70, 2, 
/* out0002_had-eta14-phi23 */     1, 70, 2, 
/* out0003_had-eta15-phi21 */     0, 
/* out0004_had-eta15-phi22 */     1, 69, 2, 
/* out0005_had-eta15-phi23 */     1, 69, 2, 
/* out0006_had-eta15-phi24 */     0, 
/* out0007_had-eta16-phi22 */     1, 69, 2, 
/* out0008_had-eta11-phi22 */     1, 71, 2, 
/* out0009_had-eta11-phi23 */     1, 71, 2, 
/* out0010_had-eta11-phi24 */     0, 
/* out0011_had-eta12-phi22 */     1, 70, 2, 
/* out0012_had-eta12-phi23 */     1, 70, 2, 
/* out0013_had-eta12-phi24 */     0, 
/* out0014_had-eta13-phi22 */     1, 70, 2, 
/* out0015_had-eta13-phi23 */     1, 70, 2, 
/* out0016_had-eta8-phi22 */     2, 83, 2, 114, 4, 
/* out0017_had-eta8-phi23 */     0, 
/* out0018_had-eta9-phi22 */     3, 71, 2, 83, 2, 114, 2, 
/* out0019_had-eta9-phi23 */     1, 71, 2, 
/* out0020_had-eta9-phi24 */     0, 
/* out0021_had-eta10-phi22 */     2, 71, 2, 113, 2, 
/* out0022_had-eta10-phi23 */     1, 71, 4, 
/* out0023_had-eta6-phi22 */     1, 106, 2, 
/* out0024_had-eta6-phi23 */     1, 106, 2, 
/* out0025_had-eta6-phi24 */     0, 
/* out0026_had-eta7-phi22 */     2, 106, 6, 115, 10, 
/* out0027_had-eta7-phi23 */     1, 106, 6, 
/* out0028_had-eta7-phi24 */     0, 
/* out0029_had-eta4-phi22 */     0, 
/* out0030_had-eta4-phi23 */     0, 
/* out0031_had-eta5-phi22 */     0, 
/* out0032_had-eta5-phi23 */     0, 
/* out0033_had-eta5-phi24 */     0, 
/* out0034_had-eta3-phi22 */     0, 
/* out0035_had-eta3-phi23 */     0, 
/* out0036_had-eta3-phi24 */     0, 
/* out0037_had-eta1-phi23 */     0, 
/* out0038_had-eta2-phi23 */     0, 
/* out0039_had-eta2-phi24 */     0, 
/* out0040_had-eta15-phi16 */     1, 37, 2, 
/* out0041_had-eta15-phi17 */     2, 37, 2, 128, 2, 
/* out0042_had-eta15-phi18 */     4, 37, 2, 81, 2, 111, 2, 128, 2, 
/* out0043_had-eta15-phi19 */     3, 37, 2, 81, 2, 111, 2, 
/* out0044_had-eta16-phi16 */     0, 
/* out0045_had-eta16-phi17 */     0, 
/* out0046_had-eta16-phi18 */     1, 111, 2, 
/* out0047_had-eta16-phi19 */     1, 111, 2, 
/* out0048_had-eta11-phi19 */     3, 38, 2, 82, 2, 129, 4, 
/* out0049_had-eta12-phi18 */     2, 38, 2, 129, 2, 
/* out0050_had-eta12-phi19 */     4, 38, 2, 82, 2, 112, 2, 129, 4, 
/* out0051_had-eta12-phi20 */     3, 38, 2, 82, 2, 112, 2, 
/* out0052_had-eta13-phi18 */     1, 128, 2, 
/* out0053_had-eta13-phi19 */     3, 38, 2, 81, 2, 112, 2, 
/* out0054_had-eta13-phi20 */     2, 81, 2, 112, 2, 
/* out0055_had-eta14-phi19 */     4, 37, 2, 81, 2, 111, 2, 128, 2, 
/* out0056_had-eta9-phi19 */     1, 130, 4, 
/* out0057_had-eta9-phi20 */     2, 83, 2, 130, 4, 
/* out0058_had-eta9-phi21 */     3, 83, 4, 113, 2, 114, 2, 
/* out0059_had-eta10-phi19 */     3, 2, 2, 38, 2, 130, 4, 
/* out0060_had-eta10-phi20 */     3, 82, 2, 113, 4, 130, 4, 
/* out0061_had-eta10-phi21 */     3, 82, 2, 83, 2, 113, 4, 
/* out0062_had-eta11-phi20 */     5, 38, 2, 82, 2, 112, 2, 113, 2, 129, 2, 
/* out0063_had-eta7-phi20 */     0, 
/* out0064_had-eta7-phi21 */     2, 114, 2, 115, 6, 
/* out0065_had-eta8-phi20 */     1, 83, 2, 
/* out0066_had-eta8-phi21 */     2, 83, 2, 114, 6, 
/* out0067_had-eta5-phi21 */     0, 
/* out0068_had-eta6-phi21 */     0, 
/* out0069_had-eta3-phi21 */     0, 
/* out0070_had-eta4-phi21 */     0, 
/* out0071_had-eta2-phi21 */     1, 147, 3, 
/* out0072_had-eta2-phi22 */     0, 
/* out0073_had-eta1-phi22 */     0, 
/* out0074_had-eta16-phi1 */     3, 84, 2, 116, 2, 131, 2, 
/* out0075_had-eta16-phi2 */     3, 84, 2, 124, 2, 131, 2, 
/* out0076_had-eta16-phi3 */     2, 124, 2, 131, 2, 
/* out0077_had-eta16-phi4 */     1, 124, 2, 
/* out0078_had-eta17-phi1 */     1, 131, 2, 
/* out0079_had-eta17-phi2 */     1, 131, 2, 
/* out0080_had-eta17-phi3 */     2, 124, 2, 131, 2, 
/* out0081_had-eta17-phi4 */     0, 
/* out0082_had-eta16-phi7 */     3, 0, 2, 9, 2, 135, 2, 
/* out0083_had-eta16-phi8 */     2, 0, 2, 9, 2, 
/* out0084_had-eta16-phi9 */     4, 0, 2, 9, 2, 34, 2, 86, 2, 
/* out0085_had-eta16-phi10 */     3, 0, 2, 34, 2, 117, 2, 
/* out0086_had-eta17-phi6 */     2, 0, 2, 9, 2, 
/* out0087_had-eta17-phi8 */     2, 0, 2, 9, 2, 
/* out0088_had-eta17-phi9 */     2, 0, 2, 9, 2, 
/* out0089_had-eta17-phi10 */     2, 0, 2, 9, 2, 
/* out0090_had-eta14-phi12 */     1, 107, 2, 
/* out0091_had-eta14-phi13 */     0, 
/* out0092_had-eta14-phi14 */     0, 
/* out0093_had-eta15-phi12 */     1, 117, 2, 
/* out0094_had-eta15-phi13 */     0, 
/* out0095_had-eta15-phi14 */     0, 
/* out0096_had-eta16-phi12 */     0, 
/* out0097_had-eta16-phi13 */     0, 
/* out0098_had-eta12-phi15 */     2, 1, 2, 39, 2, 
/* out0099_had-eta12-phi16 */     3, 1, 2, 39, 2, 132, 4, 
/* out0100_had-eta12-phi17 */     3, 1, 2, 39, 2, 132, 2, 
/* out0101_had-eta13-phi15 */     1, 1, 2, 
/* out0102_had-eta13-phi16 */     2, 1, 2, 39, 2, 
/* out0103_had-eta13-phi17 */     3, 1, 2, 37, 2, 128, 2, 
/* out0104_had-eta14-phi15 */     1, 1, 2, 
/* out0105_had-eta14-phi16 */     2, 1, 2, 128, 2, 
/* out0106_had-eta9-phi17 */     2, 2, 2, 133, 4, 
/* out0107_had-eta9-phi18 */     2, 2, 2, 133, 4, 
/* out0108_had-eta10-phi16 */     4, 2, 2, 5, 2, 39, 2, 136, 4, 
/* out0109_had-eta10-phi17 */     2, 2, 2, 133, 4, 
/* out0110_had-eta10-phi18 */     2, 2, 2, 133, 4, 
/* out0111_had-eta11-phi17 */     3, 2, 2, 39, 2, 132, 4, 
/* out0112_had-eta11-phi18 */     3, 2, 2, 38, 2, 129, 4, 
/* out0113_had-eta7-phi18 */     1, 155, 2, 
/* out0114_had-eta7-phi19 */     1, 155, 2, 
/* out0115_had-eta8-phi18 */     1, 155, 1, 
/* out0116_had-eta8-phi19 */     1, 155, 1, 
/* out0117_had-eta5-phi19 */     3, 73, 4, 141, 4, 155, 3, 
/* out0118_had-eta5-phi20 */     0, 
/* out0119_had-eta6-phi19 */     2, 141, 3, 155, 2, 
/* out0120_had-eta6-phi20 */     0, 
/* out0121_had-eta4-phi19 */     3, 73, 8, 141, 1, 156, 1, 
/* out0122_had-eta4-phi20 */     2, 73, 2, 74, 2, 
/* out0123_had-eta2-phi20 */     1, 147, 3, 
/* out0124_had-eta3-phi20 */     1, 74, 8, 
/* out0125_had-eta1-phi20 */     1, 147, 5, 
/* out0126_had-eta1-phi21 */     1, 147, 5, 
/* out0127_had-eta0-phi21 */     1, 148, 8, 
/* out0128_had-eta0-phi22 */     0, 
/* out0129_had-eta12-phi1 */     4, 87, 2, 97, 2, 118, 2, 137, 2, 
/* out0130_had-eta12-phi2 */     3, 87, 2, 125, 2, 126, 2, 
/* out0131_had-eta13-phi1 */     4, 87, 2, 96, 2, 118, 2, 134, 2, 
/* out0132_had-eta13-phi2 */     2, 125, 2, 134, 2, 
/* out0133_had-eta13-phi3 */     1, 125, 2, 
/* out0134_had-eta14-phi1 */     4, 84, 2, 96, 2, 116, 2, 134, 2, 
/* out0135_had-eta14-phi2 */     4, 84, 2, 96, 2, 125, 2, 134, 2, 
/* out0136_had-eta14-phi3 */     2, 84, 2, 125, 2, 
/* out0137_had-eta13-phi4 */     4, 3, 2, 54, 2, 75, 2, 125, 2, 
/* out0138_had-eta13-phi5 */     4, 3, 2, 54, 2, 75, 2, 98, 2, 
/* out0139_had-eta13-phi6 */     4, 3, 2, 56, 2, 88, 2, 98, 2, 
/* out0140_had-eta13-phi7 */     5, 3, 2, 56, 2, 88, 2, 93, 2, 135, 2, 
/* out0141_had-eta14-phi4 */     3, 3, 2, 53, 2, 125, 2, 
/* out0142_had-eta14-phi5 */     3, 3, 2, 53, 2, 85, 2, 
/* out0143_had-eta14-phi6 */     6, 3, 2, 53, 2, 56, 2, 85, 2, 93, 2, 135, 2, 
/* out0144_had-eta14-phi7 */     6, 3, 2, 53, 2, 56, 2, 88, 2, 93, 2, 135, 2, 
/* out0145_had-eta12-phi9 */     8, 4, 2, 10, 2, 35, 2, 58, 2, 76, 2, 89, 2, 94, 2, 138, 2, 
/* out0146_had-eta12-phi10 */     6, 4, 2, 35, 2, 76, 2, 89, 2, 108, 2, 119, 2, 
/* out0147_had-eta13-phi8 */     6, 4, 2, 10, 2, 56, 2, 88, 2, 93, 2, 138, 2, 
/* out0148_had-eta13-phi9 */     3, 4, 2, 10, 2, 72, 2, 
/* out0149_had-eta13-phi10 */     6, 4, 2, 10, 2, 35, 2, 72, 2, 89, 2, 107, 2, 
/* out0150_had-eta14-phi8 */     7, 4, 2, 10, 2, 56, 2, 72, 2, 86, 2, 93, 2, 135, 2, 
/* out0151_had-eta14-phi9 */     5, 4, 2, 10, 2, 72, 2, 86, 2, 107, 2, 
/* out0152_had-eta14-phi10 */     7, 4, 2, 10, 2, 34, 2, 72, 2, 86, 2, 107, 2, 117, 2, 
/* out0153_had-eta11-phi12 */     1, 108, 2, 
/* out0154_had-eta11-phi13 */     0, 
/* out0155_had-eta12-phi11 */     5, 35, 2, 76, 2, 89, 2, 108, 2, 119, 4, 
/* out0156_had-eta12-phi12 */     3, 35, 2, 108, 2, 119, 2, 
/* out0157_had-eta12-phi13 */     0, 
/* out0158_had-eta12-phi14 */     0, 
/* out0159_had-eta13-phi12 */     0, 
/* out0160_had-eta13-phi13 */     0, 
/* out0161_had-eta9-phi14 */     1, 5, 2, 
/* out0162_had-eta9-phi15 */     2, 5, 2, 136, 4, 
/* out0163_had-eta9-phi16 */     2, 5, 2, 136, 4, 
/* out0164_had-eta10-phi14 */     1, 5, 2, 
/* out0165_had-eta10-phi15 */     2, 5, 2, 136, 4, 
/* out0166_had-eta11-phi14 */     1, 5, 2, 
/* out0167_had-eta11-phi15 */     3, 5, 2, 39, 2, 132, 2, 
/* out0168_had-eta7-phi16 */     0, 
/* out0169_had-eta7-phi17 */     0, 
/* out0170_had-eta8-phi15 */     0, 
/* out0171_had-eta8-phi16 */     0, 
/* out0172_had-eta8-phi17 */     0, 
/* out0173_had-eta5-phi17 */     1, 13, 6, 
/* out0174_had-eta5-phi18 */     2, 141, 4, 155, 3, 
/* out0175_had-eta6-phi17 */     0, 
/* out0176_had-eta6-phi18 */     2, 141, 3, 155, 2, 
/* out0177_had-eta4-phi18 */     4, 73, 2, 77, 2, 141, 1, 156, 1, 
/* out0178_had-eta2-phi19 */     2, 142, 1, 156, 1, 
/* out0179_had-eta3-phi18 */     3, 77, 10, 142, 1, 156, 1, 
/* out0180_had-eta3-phi19 */     4, 74, 6, 77, 4, 142, 1, 156, 1, 
/* out0181_had-eta1-phi19 */     2, 142, 2, 156, 1, 
/* out0182_had-eta0-phi20 */     1, 148, 8, 
/* out0183_had-eta9-phi1 */     5, 90, 4, 99, 2, 120, 2, 127, 6, 139, 6, 
/* out0184_had-eta9-phi2 */     4, 55, 2, 78, 2, 90, 2, 127, 8, 
/* out0185_had-eta10-phi0 */     5, 90, 2, 97, 2, 99, 2, 120, 4, 139, 2, 
/* out0186_had-eta10-phi1 */     5, 90, 2, 97, 2, 120, 2, 137, 2, 139, 4, 
/* out0187_had-eta10-phi2 */     4, 55, 2, 78, 2, 126, 4, 127, 2, 
/* out0188_had-eta11-phi0 */     4, 87, 2, 97, 2, 118, 4, 137, 4, 
/* out0189_had-eta11-phi1 */     5, 87, 4, 97, 4, 118, 2, 126, 2, 137, 4, 
/* out0190_had-eta11-phi2 */     3, 87, 2, 126, 4, 137, 2, 
/* out0191_had-eta10-phi3 */     4, 6, 2, 55, 2, 78, 4, 126, 2, 
/* out0192_had-eta10-phi4 */     4, 6, 2, 55, 2, 78, 2, 100, 4, 
/* out0193_had-eta10-phi5 */     4, 6, 2, 14, 2, 57, 2, 100, 4, 
/* out0194_had-eta11-phi3 */     4, 6, 2, 54, 2, 75, 2, 126, 2, 
/* out0195_had-eta11-phi4 */     5, 6, 2, 54, 2, 57, 2, 75, 2, 100, 2, 
/* out0196_had-eta11-phi5 */     6, 6, 2, 54, 2, 57, 2, 75, 2, 98, 2, 100, 2, 
/* out0197_had-eta12-phi4 */     4, 6, 2, 54, 2, 75, 2, 98, 2, 
/* out0198_had-eta12-phi5 */     5, 6, 2, 54, 2, 57, 2, 75, 2, 98, 2, 
/* out0199_had-eta10-phi6 */     3, 7, 2, 14, 2, 57, 2, 
/* out0200_had-eta10-phi7 */     3, 7, 2, 11, 2, 91, 2, 
/* out0201_had-eta10-phi8 */     7, 7, 2, 11, 2, 58, 4, 91, 4, 94, 2, 95, 2, 140, 4, 
/* out0202_had-eta11-phi6 */     4, 7, 2, 11, 2, 57, 2, 98, 2, 
/* out0203_had-eta11-phi7 */     7, 7, 2, 11, 2, 57, 2, 58, 2, 88, 2, 94, 2, 138, 2, 
/* out0204_had-eta11-phi8 */     6, 7, 2, 11, 2, 58, 2, 91, 2, 94, 4, 138, 2, 
/* out0205_had-eta12-phi7 */     6, 7, 2, 11, 2, 88, 2, 94, 2, 98, 2, 138, 2, 
/* out0206_had-eta12-phi8 */     6, 7, 2, 11, 2, 58, 2, 88, 2, 94, 2, 138, 4, 
/* out0207_had-eta9-phi9 */     8, 8, 2, 15, 2, 40, 2, 79, 2, 91, 2, 92, 2, 95, 4, 140, 4, 
/* out0208_had-eta9-phi10 */     8, 8, 2, 12, 2, 36, 4, 79, 4, 92, 4, 95, 2, 109, 4, 121, 2, 
/* out0209_had-eta10-phi9 */     7, 8, 2, 12, 2, 58, 2, 76, 2, 91, 2, 95, 2, 140, 4, 
/* out0210_had-eta10-phi10 */     8, 8, 2, 12, 4, 36, 2, 76, 2, 79, 2, 92, 2, 109, 2, 121, 2, 
/* out0211_had-eta10-phi11 */     7, 8, 2, 12, 2, 36, 2, 92, 2, 108, 2, 109, 2, 121, 4, 
/* out0212_had-eta11-phi9 */     8, 8, 2, 12, 2, 58, 2, 76, 2, 89, 2, 94, 2, 138, 2, 140, 2, 
/* out0213_had-eta11-phi10 */     7, 8, 2, 12, 2, 35, 2, 76, 2, 89, 4, 108, 2, 119, 2, 
/* out0214_had-eta11-phi11 */     7, 8, 2, 12, 2, 35, 2, 76, 2, 89, 2, 108, 4, 119, 4, 
/* out0215_had-eta8-phi12 */     1, 123, 2, 
/* out0216_had-eta8-phi13 */     0, 
/* out0217_had-eta9-phi11 */     5, 36, 4, 79, 2, 92, 4, 109, 4, 121, 4, 
/* out0218_had-eta9-phi12 */     3, 36, 2, 109, 2, 121, 2, 
/* out0219_had-eta9-phi13 */     0, 
/* out0220_had-eta10-phi12 */     1, 121, 2, 
/* out0221_had-eta7-phi13 */     0, 
/* out0222_had-eta7-phi14 */     0, 
/* out0223_had-eta7-phi15 */     0, 
/* out0224_had-eta8-phi14 */     0, 
/* out0225_had-eta5-phi15 */     0, 
/* out0226_had-eta5-phi16 */     1, 13, 4, 
/* out0227_had-eta6-phi15 */     0, 
/* out0228_had-eta6-phi16 */     0, 
/* out0229_had-eta4-phi16 */     2, 13, 2, 16, 4, 
/* out0230_had-eta4-phi17 */     1, 13, 4, 
/* out0231_had-eta3-phi17 */     1, 16, 2, 
/* out0232_had-eta1-phi18 */     2, 142, 2, 156, 1, 
/* out0233_had-eta2-phi18 */     2, 142, 1, 156, 1, 
/* out0234_had-eta0-phi19 */     2, 142, 2, 156, 2, 
/* out0235_had-eta7-phi0 */     2, 101, 6, 122, 4, 
/* out0236_had-eta7-phi1 */     2, 101, 2, 122, 2, 
/* out0237_had-eta7-phi2 */     3, 17, 4, 80, 4, 104, 2, 
/* out0238_had-eta8-phi0 */     3, 99, 4, 101, 2, 122, 6, 
/* out0239_had-eta8-phi1 */     3, 90, 2, 99, 2, 122, 2, 
/* out0240_had-eta8-phi2 */     1, 80, 4, 
/* out0241_had-eta7-phi3 */     4, 17, 4, 80, 4, 102, 2, 104, 4, 
/* out0242_had-eta8-phi3 */     3, 55, 2, 80, 4, 102, 4, 
/* out0243_had-eta8-phi4 */     2, 18, 2, 102, 4, 
/* out0244_had-eta9-phi3 */     3, 55, 4, 78, 4, 102, 2, 
/* out0245_had-eta9-phi4 */     5, 14, 2, 55, 2, 78, 2, 100, 2, 102, 2, 
/* out0246_had-eta8-phi5 */     2, 14, 2, 18, 2, 
/* out0247_had-eta8-phi6 */     1, 14, 2, 
/* out0248_had-eta9-phi5 */     2, 14, 2, 100, 2, 
/* out0249_had-eta9-phi6 */     1, 14, 4, 
/* out0250_had-eta7-phi8 */     0, 
/* out0251_had-eta8-phi7 */     1, 15, 2, 
/* out0252_had-eta8-phi8 */     2, 15, 4, 40, 4, 
/* out0253_had-eta8-phi9 */     3, 15, 2, 40, 4, 95, 2, 
/* out0254_had-eta9-phi7 */     2, 15, 2, 91, 2, 
/* out0255_had-eta9-phi8 */     5, 15, 4, 40, 2, 91, 2, 95, 4, 140, 2, 
/* out0256_had-eta7-phi9 */     2, 40, 2, 41, 2, 
/* out0257_had-eta7-phi10 */     2, 41, 2, 110, 2, 
/* out0258_had-eta7-phi11 */     2, 110, 8, 123, 6, 
/* out0259_had-eta8-phi10 */     4, 40, 2, 79, 4, 92, 2, 123, 2, 
/* out0260_had-eta8-phi11 */     5, 36, 2, 79, 2, 109, 2, 110, 4, 123, 6, 
/* out0261_had-eta6-phi11 */     0, 
/* out0262_had-eta6-phi12 */     1, 145, 1, 
/* out0263_had-eta6-phi13 */     1, 145, 1, 
/* out0264_had-eta7-phi12 */     1, 110, 2, 
/* out0265_had-eta5-phi13 */     1, 145, 3, 
/* out0266_had-eta5-phi14 */     0, 
/* out0267_had-eta6-phi14 */     0, 
/* out0268_had-eta4-phi14 */     1, 149, 6, 
/* out0269_had-eta4-phi15 */     1, 149, 6, 
/* out0270_had-eta2-phi16 */     1, 19, 6, 
/* out0271_had-eta3-phi15 */     3, 16, 2, 19, 2, 149, 2, 
/* out0272_had-eta3-phi16 */     1, 16, 8, 
/* out0273_had-eta1-phi17 */     0, 
/* out0274_had-eta2-phi17 */     0, 
/* out0275_had-eta5-phi0 */     1, 103, 8, 
/* out0276_had-eta5-phi1 */     2, 20, 2, 103, 2, 
/* out0277_had-eta6-phi0 */     2, 101, 4, 103, 4, 
/* out0278_had-eta6-phi1 */     0, 
/* out0279_had-eta5-phi2 */     2, 20, 6, 105, 6, 
/* out0280_had-eta6-phi2 */     3, 17, 4, 20, 2, 104, 2, 
/* out0281_had-eta6-phi3 */     3, 17, 4, 21, 2, 104, 6, 
/* out0282_had-eta6-phi4 */     5, 18, 2, 21, 2, 59, 4, 104, 2, 151, 1, 
/* out0283_had-eta6-phi5 */     4, 18, 2, 22, 2, 59, 4, 151, 1, 
/* out0284_had-eta7-phi4 */     2, 18, 4, 102, 2, 
/* out0285_had-eta7-phi5 */     1, 18, 4, 
/* out0286_had-eta6-phi6 */     2, 22, 4, 42, 4, 
/* out0287_had-eta6-phi7 */     1, 42, 2, 
/* out0288_had-eta7-phi6 */     0, 
/* out0289_had-eta7-phi7 */     0, 
/* out0290_had-eta5-phi8 */     0, 
/* out0291_had-eta5-phi9 */     2, 41, 2, 43, 4, 
/* out0292_had-eta6-phi8 */     0, 
/* out0293_had-eta6-phi9 */     1, 41, 6, 
/* out0294_had-eta5-phi10 */     1, 43, 4, 
/* out0295_had-eta5-phi11 */     0, 
/* out0296_had-eta6-phi10 */     1, 41, 4, 
/* out0297_had-eta4-phi12 */     1, 145, 4, 
/* out0298_had-eta4-phi13 */     1, 145, 4, 
/* out0299_had-eta5-phi12 */     1, 145, 3, 
/* out0300_had-eta3-phi13 */     1, 146, 1, 
/* out0301_had-eta3-phi14 */     1, 149, 2, 
/* out0302_had-eta2-phi14 */     2, 143, 5, 150, 1, 
/* out0303_had-eta2-phi15 */     3, 19, 8, 143, 5, 150, 1, 
/* out0304_had-eta1-phi15 */     4, 23, 14, 143, 3, 144, 1, 150, 2, 
/* out0305_had-eta1-phi16 */     1, 23, 2, 
/* out0306_had-eta0-phi16 */     0, 
/* out0307_had-eta3-phi0 */     0, 
/* out0308_had-eta3-phi1 */     1, 24, 4, 
/* out0309_had-eta4-phi0 */     0, 
/* out0310_had-eta4-phi1 */     1, 24, 2, 
/* out0311_had-eta4-phi2 */     3, 20, 4, 24, 4, 105, 2, 
/* out0312_had-eta4-phi3 */     3, 25, 6, 60, 2, 105, 2, 
/* out0313_had-eta4-phi4 */     6, 21, 2, 25, 2, 26, 4, 60, 10, 151, 4, 159, 6, 
/* out0314_had-eta5-phi3 */     3, 20, 2, 21, 4, 105, 6, 
/* out0315_had-eta5-phi4 */     4, 21, 6, 59, 4, 60, 2, 151, 3, 
/* out0316_had-eta4-phi5 */     5, 26, 8, 44, 6, 60, 2, 151, 4, 159, 6, 
/* out0317_had-eta4-phi6 */     2, 44, 6, 45, 2, 
/* out0318_had-eta5-phi5 */     3, 22, 4, 59, 4, 151, 3, 
/* out0319_had-eta5-phi6 */     2, 22, 6, 42, 6, 
/* out0320_had-eta4-phi7 */     1, 45, 8, 
/* out0321_had-eta4-phi8 */     1, 45, 2, 
/* out0322_had-eta5-phi7 */     1, 42, 4, 
/* out0323_had-eta4-phi9 */     1, 43, 4, 
/* out0324_had-eta4-phi10 */     2, 43, 4, 46, 2, 
/* out0325_had-eta3-phi10 */     1, 46, 10, 
/* out0326_had-eta3-phi11 */     0, 
/* out0327_had-eta4-phi11 */     0, 
/* out0328_had-eta3-phi12 */     1, 146, 1, 
/* out0329_had-eta2-phi13 */     1, 146, 1, 
/* out0330_had-eta1-phi14 */     3, 143, 3, 144, 1, 150, 2, 
/* out0331_had-eta0-phi15 */     2, 144, 5, 150, 2, 
/* out0332_had-eta2-phi0 */     1, 153, 5, 
/* out0333_had-eta2-phi1 */     3, 27, 8, 62, 2, 153, 5, 
/* out0334_had-eta2-phi2 */     3, 27, 6, 28, 4, 31, 2, 
/* out0335_had-eta3-phi2 */     2, 24, 6, 28, 2, 
/* out0336_had-eta3-phi3 */     3, 25, 6, 28, 4, 61, 6, 
/* out0337_had-eta3-phi4 */     6, 25, 2, 26, 2, 29, 6, 61, 6, 152, 1, 159, 2, 
/* out0338_had-eta3-phi5 */     5, 26, 2, 29, 2, 44, 2, 152, 1, 159, 2, 
/* out0339_had-eta3-phi6 */     1, 44, 2, 
/* out0340_had-eta3-phi7 */     2, 45, 4, 47, 4, 
/* out0341_had-eta3-phi8 */     1, 47, 4, 
/* out0342_had-eta2-phi9 */     0, 
/* out0343_had-eta3-phi9 */     1, 46, 4, 
/* out0344_had-eta2-phi10 */     2, 48, 12, 157, 3, 
/* out0345_had-eta2-phi11 */     2, 48, 2, 157, 3, 
/* out0346_had-eta1-phi12 */     1, 146, 1, 
/* out0347_had-eta2-phi12 */     1, 146, 1, 
/* out0348_had-eta1-phi13 */     1, 146, 1, 
/* out0349_had-eta0-phi13 */     1, 146, 2, 
/* out0350_had-eta0-phi14 */     2, 144, 5, 150, 2, 
/* out0351_had-eta1-phi0 */     3, 62, 2, 153, 3, 154, 1, 
/* out0352_had-eta1-phi1 */     6, 27, 2, 30, 10, 62, 12, 66, 2, 153, 3, 154, 1, 
/* out0353_had-eta1-phi2 */     3, 30, 4, 31, 8, 66, 4, 
/* out0354_had-eta2-phi3 */     4, 28, 6, 32, 2, 61, 2, 63, 10, 
/* out0355_had-eta2-phi4 */     7, 29, 6, 32, 4, 49, 6, 61, 2, 63, 2, 152, 1, 160, 1, 
/* out0356_had-eta2-phi5 */     4, 29, 2, 49, 2, 152, 1, 160, 1, 
/* out0357_had-eta2-phi6 */     0, 
/* out0358_had-eta2-phi7 */     1, 47, 4, 
/* out0359_had-eta2-phi8 */     2, 47, 4, 50, 6, 
/* out0360_had-eta1-phi9 */     1, 67, 4, 
/* out0361_had-eta1-phi10 */     5, 48, 2, 51, 10, 64, 12, 67, 2, 157, 5, 
/* out0362_had-eta1-phi11 */     3, 51, 2, 64, 4, 157, 5, 
/* out0363_had-eta0-phi1 */     4, 30, 2, 65, 12, 66, 4, 154, 5, 
/* out0364_had-eta0-phi2 */     1, 66, 6, 
/* out0365_had-eta1-phi3 */     5, 31, 6, 32, 4, 33, 6, 52, 2, 63, 4, 
/* out0366_had-eta1-phi4 */     6, 32, 6, 33, 2, 49, 6, 52, 8, 152, 1, 160, 2, 
/* out0367_had-eta1-phi5 */     3, 49, 2, 152, 1, 160, 2, 
/* out0368_had-eta1-phi6 */     0, 
/* out0369_had-eta1-phi7 */     1, 50, 2, 
/* out0370_had-eta1-phi8 */     1, 50, 8, 
/* out0371_had-eta0-phi9 */     1, 67, 6, 
/* out0372_had-eta0-phi10 */     4, 51, 4, 67, 4, 68, 12, 158, 8, 
/* out0373_had-eta16-phi20 */     1, 111, 2, 
/* out0374_had-eta16-phi21 */     1, 69, 2, 
/* out0375_had-eta17-phi19 */     0, 
/* out0376_had-eta17-phi20 */     0, 
/* out0377_had-eta17-phi21 */     1, 69, 2, 
/* out0378_had-eta17-phi22 */     1, 69, 2, 
/* out0379_had-eta12-phi21 */     2, 82, 2, 112, 4, 
/* out0380_had-eta13-phi21 */     2, 70, 2, 112, 2, 
/* out0381_had-eta14-phi20 */     2, 81, 2, 111, 2, 
/* out0382_had-eta11-phi21 */     2, 82, 2, 113, 2, 
/* out0383_had-eta16-phi14 */     0, 
/* out0384_had-eta16-phi15 */     0, 
/* out0385_had-eta17-phi13 */     0, 
/* out0386_had-eta17-phi14 */     0, 
/* out0387_had-eta17-phi15 */     0, 
/* out0388_had-eta17-phi16 */     0, 
/* out0389_had-eta17-phi17 */     0, 
/* out0390_had-eta14-phi17 */     2, 37, 2, 128, 2, 
/* out0391_had-eta14-phi18 */     3, 37, 2, 81, 2, 128, 2, 
/* out0392_had-eta14-phi0 */     3, 96, 2, 116, 2, 134, 2, 
/* out0393_had-eta15-phi0 */     2, 96, 2, 116, 2, 
/* out0394_had-eta15-phi1 */     4, 84, 2, 96, 2, 116, 2, 134, 2, 
/* out0395_had-eta15-phi2 */     4, 84, 2, 116, 2, 131, 2, 134, 2, 
/* out0396_had-eta16-phi0 */     2, 116, 2, 131, 2, 
/* out0397_had-eta15-phi4 */     3, 53, 2, 85, 2, 124, 2, 
/* out0398_had-eta15-phi5 */     3, 53, 2, 85, 2, 124, 2, 
/* out0399_had-eta15-phi6 */     4, 53, 2, 85, 2, 93, 2, 135, 2, 
/* out0400_had-eta16-phi5 */     2, 85, 2, 124, 2, 
/* out0401_had-eta16-phi6 */     1, 85, 2, 
/* out0402_had-eta14-phi11 */     2, 107, 2, 117, 2, 
/* out0403_had-eta15-phi9 */     5, 10, 2, 34, 2, 72, 2, 86, 2, 117, 2, 
/* out0404_had-eta15-phi10 */     5, 34, 2, 72, 2, 86, 2, 107, 2, 117, 2, 
/* out0405_had-eta15-phi11 */     4, 34, 2, 86, 2, 107, 2, 117, 2, 
/* out0406_had-eta16-phi11 */     2, 34, 2, 117, 2, 
/* out0407_had-eta13-phi14 */     0, 
/* out0408_had-eta11-phi16 */     2, 39, 2, 132, 4, 
/* out0409_had-eta12-phi-1 */     1, 118, 2, 
/* out0410_had-eta12-phi0 */     4, 87, 2, 97, 2, 118, 2, 137, 2, 
/* out0411_had-eta13-phi0 */     3, 96, 2, 118, 2, 134, 2, 
/* out0412_had-eta12-phi3 */     3, 54, 2, 75, 2, 125, 2, 
/* out0413_had-eta12-phi6 */     4, 11, 2, 57, 2, 88, 2, 98, 2, 
/* out0414_had-eta13-phi11 */     3, 35, 2, 107, 2, 119, 2, 
/* out0415_had-eta10-phi13 */     0, 
/* out0416_had-eta9-phi-1 */     2, 99, 2, 120, 2, 
/* out0417_had-eta9-phi0 */     4, 90, 4, 99, 4, 120, 4, 139, 4, 
/* out0418_had-eta0-phi18 */     2, 142, 2, 156, 2, 
/* out0419_had-eta7-phi-1 */     1, 101, 2, 
/* out0420_had-eta5-phi-1 */     1, 103, 2, 
/* out0421_had-eta0-phi17 */     0, 
/* out0422_had-eta3-phi-1 */     0, 
/* out0423_had-eta2-phi-1 */     0, 
/* out0424_had-eta0-phi0 */     2, 65, 4, 154, 5, 
/* out0425_had-eta1-phi-1 */     0, 
/* out0426_had-eta0-phi11 */     2, 68, 4, 158, 8, 
/* out0427_had-eta0-phi3 */     2, 33, 6, 52, 2, 
/* out0428_had-eta0-phi8 */     0, 
/* out0429_had-eta16-phi23 */     1, 69, 2, 
/* out0430_had-eta4-phi24 */     0, 
/* out0431_had-eta0-phi23 */     0, 
/* out0432_had-eta1-phi24 */     0, 
/* out0433_had-eta17-phi5 */     0, 
/* out0434_had-eta17-phi7 */     1, 9, 2, 
/* out0435_had-eta0-phi12 */     1, 146, 2, 
/* out0436_had-eta0-phi4 */     4, 33, 2, 52, 4, 152, 2, 160, 2, 
/* out0437_had-eta0-phi5 */     2, 152, 2, 160, 2, 
/* out0438_had-eta0-phi6 */     0, 
/* out0439_had-eta0-phi7 */     0, 
/* out0440_had-eta17-phi18 */     0, 
/* out0441_had-eta16-phi-1 */     0, 
/* out0442_had-eta17-phi11 */     1, 34, 2, 
/* out0443_had-eta4-phi-1 */     0, 
/* out0444_had-eta16-phi24 */     0, 
/* out0445_had-eta17-phi23 */     1, 69, 2, 
/* out0446_had-eta10-phi24 */     1, 71, 2, 
/* out0447_had-eta17-phi12 */     0, 
/* out0448_had-eta15-phi7 */     5, 53, 2, 56, 2, 85, 2, 93, 2, 135, 2, 
/* out0449_had-eta17-phi0 */     0, 
/* out0450_had-eta15-phi15 */     0, 
/* out0451_had-eta10-phi-1 */     1, 120, 2, 
/* out0452_had-eta8-phi-1 */     1, 122, 2, 
/* out0453_had-eta13-phi24 */     1, 70, 2, 
/* out0454_had-eta8-phi24 */     0, 
/* out0455_had-eta0-phi24 */     0, 
/* out0456_had-eta15-phi8 */     5, 56, 2, 72, 2, 86, 2, 93, 2, 135, 2, 
/* out0457_had-eta13-phi-1 */     0, 
/* out0458_had-eta15-phi3 */     2, 84, 2, 124, 2, 
/* out0459_had-eta6-phi-1 */     0, 
/* out0460_had-eta15-phi20 */     2, 81, 2, 111, 2, 
/* out0461_had-eta17-phi24 */     0, 
/* out0462_had-eta17-phi-1 */     0, 
/* out0463_had-eta11-phi-1 */     1, 97, 2, 
/* out0464_had-eta14-phi24 */     0, 
/* out0465_had-eta14-phi-1 */     1, 96, 2, 
/* out0466_had-eta15-phi-1 */     1, 116, 2, 
/* out0467_had-eta-2-phi0 */     0, 
/* out0468_had-eta-1-phi0 */     1, 154, 2, 
/* out0469_had-eta-2-phi1 */     0, 
/* out0470_had-eta-1-phi1 */     1, 154, 2, 
/* out0471_had-eta-2-phi2 */     0, 
/* out0472_had-eta-1-phi2 */     0, 
/* out0473_had-eta-2-phi3 */     0, 
/* out0474_had-eta-1-phi3 */     0, 
/* out0475_had-eta-2-phi4 */     1, 152, 1, 
/* out0476_had-eta-1-phi4 */     2, 152, 2, 160, 3, 
/* out0477_had-eta-2-phi5 */     1, 152, 1, 
/* out0478_had-eta-1-phi5 */     2, 152, 2, 160, 3, 
/* out0479_had-eta-2-phi6 */     0, 
/* out0480_had-eta-1-phi6 */     0, 
/* out0481_had-eta-2-phi7 */     0, 
/* out0482_had-eta-1-phi7 */     0, 
/* out0483_had-eta-2-phi8 */     0, 
/* out0484_had-eta-1-phi8 */     0, 
/* out0485_had-eta-2-phi9 */     0, 
/* out0486_had-eta-1-phi9 */     0, 
/* out0487_had-eta-2-phi10 */     0, 
/* out0488_had-eta-1-phi10 */     0, 
/* out0489_had-eta-2-phi11 */     0, 
/* out0490_had-eta-1-phi11 */     0, 
/* out0491_had-eta-2-phi12 */     1, 146, 1, 
/* out0492_had-eta-1-phi12 */     1, 146, 2, 
/* out0493_had-eta-2-phi13 */     1, 146, 1, 
/* out0494_had-eta-1-phi13 */     1, 146, 2, 
/* out0495_had-eta-2-phi14 */     0, 
/* out0496_had-eta-1-phi14 */     2, 144, 2, 150, 3, 
/* out0497_had-eta-2-phi15 */     0, 
/* out0498_had-eta-1-phi15 */     2, 144, 2, 150, 3, 
/* out0499_had-eta-2-phi16 */     0, 
/* out0500_had-eta-1-phi16 */     0, 
/* out0501_had-eta-2-phi17 */     0, 
/* out0502_had-eta-1-phi17 */     0, 
/* out0503_had-eta-2-phi18 */     0, 
/* out0504_had-eta-1-phi18 */     2, 142, 2, 156, 2, 
/* out0505_had-eta-2-phi19 */     0, 
/* out0506_had-eta-1-phi19 */     2, 142, 2, 156, 2, 
/* out0507_had-eta-2-phi20 */     0, 
/* out0508_had-eta-1-phi20 */     0, 
/* out0509_had-eta-2-phi21 */     0, 
/* out0510_had-eta-1-phi21 */     0, 
/* out0511_had-eta-2-phi22 */     0, 
/* out0512_had-eta-1-phi22 */     0, 
/* out0513_had-eta-2-phi23 */     0, 
/* out0514_had-eta-1-phi23 */     0
};